`timescale 1ns / 1ps
module non_restoring_division(
	input [31:0] M,
	input [31:0] D,
	output [31:0] R,
	output [31:0] Q
	);
// Level - 1
	wire [3:0] OUT_0_0;
	CAS CAS_0_0( {1'b1, D[31], M[0], 1'b1}, OUT_0_0);
	wire [3:0] OUT_0_1;
	CAS CAS_0_1( { OUT_0_0[0], 1'b0, M[1], 1'b1}, OUT_0_1);
        wire [3:0] OUT_0_2;
        CAS CAS_0_2( { OUT_0_1[0], 1'b0, M[2], 1'b1}, OUT_0_2);
        wire [3:0] OUT_0_3;
        CAS CAS_0_3( { OUT_0_2[0], 1'b0, M[3], 1'b1}, OUT_0_3);
        wire [3:0] OUT_0_4;
        CAS CAS_0_4( { OUT_0_3[0], 1'b0, M[4], 1'b1}, OUT_0_4);
        wire [3:0] OUT_0_5;
        CAS CAS_0_5( { OUT_0_4[0], 1'b0, M[5], 1'b1}, OUT_0_5);
        wire [3:0] OUT_0_6;
        CAS CAS_0_6( { OUT_0_5[0], 1'b0, M[6], 1'b1}, OUT_0_6);
        wire [3:0] OUT_0_7;
        CAS CAS_0_7( { OUT_0_6[0], 1'b0, M[7], 1'b1}, OUT_0_7);
        wire [3:0] OUT_0_8;
        CAS CAS_0_8( { OUT_0_7[0], 1'b0, M[8], 1'b1}, OUT_0_8);
        wire [3:0] OUT_0_9;
        CAS CAS_0_9( { OUT_0_8[0], 1'b0, M[9], 1'b1}, OUT_0_9);
        wire [3:0] OUT_0_10;
        CAS CAS_0_10( { OUT_0_9[0], 1'b0, M[10], 1'b1}, OUT_0_10);
        wire [3:0] OUT_0_11;
        CAS CAS_0_11( { OUT_0_10[0], 1'b0, M[11], 1'b1}, OUT_0_11);
        wire [3:0] OUT_0_12;
        CAS CAS_0_12( { OUT_0_11[0], 1'b0, M[12], 1'b1}, OUT_0_12);
        wire [3:0] OUT_0_13;
        CAS CAS_0_13( { OUT_0_12[0], 1'b0, M[13], 1'b1}, OUT_0_13);
        wire [3:0] OUT_0_14;
        CAS CAS_0_14( { OUT_0_13[0], 1'b0, M[14], 1'b1}, OUT_0_14);
        wire [3:0] OUT_0_15;
        CAS CAS_0_15( { OUT_0_14[0], 1'b0, M[15], 1'b1}, OUT_0_15);
        wire [3:0] OUT_0_16;
        CAS CAS_0_16( { OUT_0_15[0], 1'b0, M[16], 1'b1}, OUT_0_16);
        wire [3:0] OUT_0_17;
        CAS CAS_0_17( { OUT_0_16[0], 1'b0, M[17], 1'b1}, OUT_0_17);
        wire [3:0] OUT_0_18;
        CAS CAS_0_18( { OUT_0_17[0], 1'b0, M[18], 1'b1}, OUT_0_18);
        wire [3:0] OUT_0_19;
        CAS CAS_0_19( { OUT_0_18[0], 1'b0, M[19], 1'b1}, OUT_0_19);
        wire [3:0] OUT_0_20;
        CAS CAS_0_20( { OUT_0_19[0], 1'b0, M[20], 1'b1}, OUT_0_20);
        wire [3:0] OUT_0_21;
        CAS CAS_0_21( { OUT_0_20[0], 1'b0, M[21], 1'b1}, OUT_0_21);
        wire [3:0] OUT_0_22;
        CAS CAS_0_22( { OUT_0_21[0], 1'b0, M[22], 1'b1}, OUT_0_22);
        wire [3:0] OUT_0_23;
        CAS CAS_0_23( { OUT_0_22[0], 1'b0, M[23], 1'b1}, OUT_0_23);
        wire [3:0] OUT_0_24;
        CAS CAS_0_24( { OUT_0_23[0], 1'b0, M[24], 1'b1}, OUT_0_24);
        wire [3:0] OUT_0_25;
        CAS CAS_0_25( { OUT_0_24[0], 1'b0, M[25], 1'b1}, OUT_0_25);
        wire [3:0] OUT_0_26;
        CAS CAS_0_26( { OUT_0_25[0], 1'b0, M[26], 1'b1}, OUT_0_26);
        wire [3:0] OUT_0_27;
        CAS CAS_0_27( { OUT_0_26[0], 1'b0, M[27], 1'b1}, OUT_0_27);
        wire [3:0] OUT_0_28;
        CAS CAS_0_28( { OUT_0_27[0], 1'b0, M[28], 1'b1}, OUT_0_28);
        wire [3:0] OUT_0_29;
        CAS CAS_0_29( { OUT_0_28[0], 1'b0, M[29], 1'b1}, OUT_0_29);
        wire [3:0] OUT_0_30;
        CAS CAS_0_30( { OUT_0_29[0], 1'b0, M[30], 1'b1}, OUT_0_30);
        wire [3:0] OUT_0_31;
        CAS CAS_0_31( { OUT_0_30[0], 1'b0, M[31], 1'b1}, OUT_0_31);
	assign Q[31] = OUT_0_31[0];

// Level - 2
	wire [3:0] OUT_1_0;
        CAS CAS_1_0( {Q[31], D[30], M[0], Q[31]}, OUT_1_0);
        wire [3:0] OUT_1_1;
        CAS CAS_1_1( { OUT_1_0[0], OUT_0_0[1], M[1], Q[31]}, OUT_1_1);
        wire [3:0] OUT_1_2;
        CAS CAS_1_2( { OUT_1_1[0], OUT_0_1[1], M[2], Q[31]}, OUT_1_2);
        wire [3:0] OUT_1_3;
        CAS CAS_1_3( { OUT_1_2[0], OUT_0_2[1], M[3], Q[31]}, OUT_1_3);
        wire [3:0] OUT_1_4;
        CAS CAS_1_4( { OUT_1_3[0], OUT_0_3[1], M[4], Q[31]}, OUT_1_4);
        wire [3:0] OUT_1_5;
        CAS CAS_1_5( { OUT_1_4[0], OUT_0_4[1], M[5], Q[31]}, OUT_1_5);
        wire [3:0] OUT_1_6;
        CAS CAS_1_6( { OUT_1_5[0], OUT_0_5[1], M[6], Q[31]}, OUT_1_6);
        wire [3:0] OUT_1_7;
        CAS CAS_1_7( { OUT_1_6[0], OUT_0_6[1], M[7], Q[31]}, OUT_1_7);
        wire [3:0] OUT_1_8;
        CAS CAS_1_8( { OUT_1_7[0], OUT_0_7[1], M[8], Q[31]}, OUT_1_8);
        wire [3:0] OUT_1_9;
        CAS CAS_1_9( { OUT_1_8[0], OUT_0_8[1], M[9], Q[31]}, OUT_1_9);
        wire [3:0] OUT_1_10;
        CAS CAS_1_10( { OUT_1_9[0], OUT_0_9[1], M[10], Q[31]}, OUT_1_10);
        wire [3:0] OUT_1_11;
        CAS CAS_1_11( { OUT_1_10[0], OUT_0_10[1], M[11], Q[31]}, OUT_1_11);
        wire [3:0] OUT_1_12;
        CAS CAS_1_12( { OUT_1_11[0], OUT_0_11[1], M[12], Q[31]}, OUT_1_12);
        wire [3:0] OUT_1_13;
        CAS CAS_1_13( { OUT_1_12[0], OUT_0_12[1], M[13], Q[31]}, OUT_1_13);
        wire [3:0] OUT_1_14;
        CAS CAS_1_14( { OUT_1_13[0], OUT_0_13[1], M[14], Q[31]}, OUT_1_14);
        wire [3:0] OUT_1_15;
        CAS CAS_1_15( { OUT_1_14[0], OUT_0_14[1], M[15], Q[31]}, OUT_1_15);
        wire [3:0] OUT_1_16;
        CAS CAS_1_16( { OUT_1_15[0], OUT_0_15[1], M[16], Q[31]}, OUT_1_16);
        wire [3:0] OUT_1_17;
        CAS CAS_1_17( { OUT_1_16[0], OUT_0_16[1], M[17], Q[31]}, OUT_1_17);
        wire [3:0] OUT_1_18;
        CAS CAS_1_18( { OUT_1_17[0], OUT_0_17[1], M[18], Q[31]}, OUT_1_18);
        wire [3:0] OUT_1_19;
        CAS CAS_1_19( { OUT_1_18[0], OUT_0_18[1], M[19], Q[31]}, OUT_1_19);
        wire [3:0] OUT_1_20;
        CAS CAS_1_20( { OUT_1_19[0], OUT_0_19[1], M[20], Q[31]}, OUT_1_20);
        wire [3:0] OUT_1_21;
        CAS CAS_1_21( { OUT_1_20[0], OUT_0_20[1], M[21], Q[31]}, OUT_1_21);
        wire [3:0] OUT_1_22;
        CAS CAS_1_22( { OUT_1_21[0], OUT_0_21[1], M[22], Q[31]}, OUT_1_22);
        wire [3:0] OUT_1_23;
        CAS CAS_1_23( { OUT_1_22[0], OUT_0_22[1], M[23], Q[31]}, OUT_1_23);
        wire [3:0] OUT_1_24;
        CAS CAS_1_24( { OUT_1_23[0], OUT_0_23[1], M[24], Q[31]}, OUT_1_24);
        wire [3:0] OUT_1_25;
        CAS CAS_1_25( { OUT_1_24[0], OUT_0_24[1], M[25], Q[31]}, OUT_1_25);
        wire [3:0] OUT_1_26;
        CAS CAS_1_26( { OUT_1_25[0], OUT_0_25[1], M[26], Q[31]}, OUT_1_26);
        wire [3:0] OUT_1_27;
        CAS CAS_1_27( { OUT_1_26[0], OUT_0_26[1], M[27], Q[31]}, OUT_1_27);
        wire [3:0] OUT_1_28;
        CAS CAS_1_28( { OUT_1_27[0], OUT_0_27[1], M[28], Q[31]}, OUT_1_28);
        wire [3:0] OUT_1_29;
        CAS CAS_1_29( { OUT_1_28[0], OUT_0_28[1], M[29], Q[31]}, OUT_1_29);
        wire [3:0] OUT_1_30;
        CAS CAS_1_30( { OUT_1_29[0], OUT_0_29[1], M[30], Q[31]}, OUT_1_30);
        wire [3:0] OUT_1_31;
        CAS CAS_1_31( { OUT_1_30[0], OUT_0_30[1], M[31], Q[31]}, OUT_1_31);
        assign Q[30] = OUT_1_31[0];

// Level - 3
	wire [3:0] OUT_2_0;
	CAS CAS_2_0( {Q[30], D[29], M[0], Q[30]}, OUT_2_0);
	wire [3:0] OUT_2_1;
	CAS CAS_2_1( {OUT_2_0[0], OUT_1_0[1], M[1], Q[30]}, OUT_2_1);
	wire [3:0] OUT_2_2;
	CAS CAS_2_2( {OUT_2_1[0], OUT_1_1[1], M[2], Q[30]}, OUT_2_2);
	wire [3:0] OUT_2_3;
	CAS CAS_2_3( {OUT_2_2[0], OUT_1_2[1], M[3], Q[30]}, OUT_2_3);
	wire [3:0] OUT_2_4;
	CAS CAS_2_4( {OUT_2_3[0], OUT_1_3[1], M[4], Q[30]}, OUT_2_4);
	wire [3:0] OUT_2_5;
	CAS CAS_2_5( {OUT_2_4[0], OUT_1_4[1], M[5], Q[30]}, OUT_2_5);
	wire [3:0] OUT_2_6;
	CAS CAS_2_6( {OUT_2_5[0], OUT_1_5[1], M[6], Q[30]}, OUT_2_6);
	wire [3:0] OUT_2_7;
	CAS CAS_2_7( {OUT_2_6[0], OUT_1_6[1], M[7], Q[30]}, OUT_2_7);
	wire [3:0] OUT_2_8;
	CAS CAS_2_8( {OUT_2_7[0], OUT_1_7[1], M[8], Q[30]}, OUT_2_8);
	wire [3:0] OUT_2_9;
	CAS CAS_2_9( {OUT_2_8[0], OUT_1_8[1], M[9], Q[30]}, OUT_2_9);
	wire [3:0] OUT_2_10;
	CAS CAS_2_10( {OUT_2_9[0], OUT_1_9[1], M[10], Q[30]}, OUT_2_10);
	wire [3:0] OUT_2_11;
	CAS CAS_2_11( {OUT_2_10[0], OUT_1_10[1], M[11], Q[30]}, OUT_2_11);
	wire [3:0] OUT_2_12;
	CAS CAS_2_12( {OUT_2_11[0], OUT_1_11[1], M[12], Q[30]}, OUT_2_12);
	wire [3:0] OUT_2_13;
	CAS CAS_2_13( {OUT_2_12[0], OUT_1_12[1], M[13], Q[30]}, OUT_2_13);
	wire [3:0] OUT_2_14;
	CAS CAS_2_14( {OUT_2_13[0], OUT_1_13[1], M[14], Q[30]}, OUT_2_14);
	wire [3:0] OUT_2_15;
	CAS CAS_2_15( {OUT_2_14[0], OUT_1_14[1], M[15], Q[30]}, OUT_2_15);
	wire [3:0] OUT_2_16;
	CAS CAS_2_16( {OUT_2_15[0], OUT_1_15[1], M[16], Q[30]}, OUT_2_16);
	wire [3:0] OUT_2_17;
	CAS CAS_2_17( {OUT_2_16[0], OUT_1_16[1], M[17], Q[30]}, OUT_2_17);
	wire [3:0] OUT_2_18;
	CAS CAS_2_18( {OUT_2_17[0], OUT_1_17[1], M[18], Q[30]}, OUT_2_18);
	wire [3:0] OUT_2_19;
	CAS CAS_2_19( {OUT_2_18[0], OUT_1_18[1], M[19], Q[30]}, OUT_2_19);
	wire [3:0] OUT_2_20;
	CAS CAS_2_20( {OUT_2_19[0], OUT_1_19[1], M[20], Q[30]}, OUT_2_20);
	wire [3:0] OUT_2_21;
	CAS CAS_2_21( {OUT_2_20[0], OUT_1_20[1], M[21], Q[30]}, OUT_2_21);
	wire [3:0] OUT_2_22;
	CAS CAS_2_22( {OUT_2_21[0], OUT_1_21[1], M[22], Q[30]}, OUT_2_22);
	wire [3:0] OUT_2_23;
	CAS CAS_2_23( {OUT_2_22[0], OUT_1_22[1], M[23], Q[30]}, OUT_2_23);
	wire [3:0] OUT_2_24;
	CAS CAS_2_24( {OUT_2_23[0], OUT_1_23[1], M[24], Q[30]}, OUT_2_24);
	wire [3:0] OUT_2_25;
	CAS CAS_2_25( {OUT_2_24[0], OUT_1_24[1], M[25], Q[30]}, OUT_2_25);
	wire [3:0] OUT_2_26;
	CAS CAS_2_26( {OUT_2_25[0], OUT_1_25[1], M[26], Q[30]}, OUT_2_26);
	wire [3:0] OUT_2_27;
	CAS CAS_2_27( {OUT_2_26[0], OUT_1_26[1], M[27], Q[30]}, OUT_2_27);
	wire [3:0] OUT_2_28;
	CAS CAS_2_28( {OUT_2_27[0], OUT_1_27[1], M[28], Q[30]}, OUT_2_28);
	wire [3:0] OUT_2_29;
	CAS CAS_2_29( {OUT_2_28[0], OUT_1_28[1], M[29], Q[30]}, OUT_2_29);
	wire [3:0] OUT_2_30;
	CAS CAS_2_30( {OUT_2_29[0], OUT_1_29[1], M[30], Q[30]}, OUT_2_30);
	wire [3:0] OUT_2_31;
	CAS CAS_2_31( {OUT_2_30[0], OUT_1_30[1], M[31], Q[30]}, OUT_2_31);
	assign Q[29] = OUT_2_31[0];

// Level - 4
	wire [3:0] OUT_3_0;
	CAS CAS_3_0( {Q[29], D[28], M[0], Q[29]}, OUT_3_0);
	wire [3:0] OUT_3_1;
	CAS CAS_3_1( {OUT_3_0[0], OUT_2_0[1], M[1], Q[29]}, OUT_3_1);
	wire [3:0] OUT_3_2;
	CAS CAS_3_2( {OUT_3_1[0], OUT_2_1[1], M[2], Q[29]}, OUT_3_2);
	wire [3:0] OUT_3_3;
	CAS CAS_3_3( {OUT_3_2[0], OUT_2_2[1], M[3], Q[29]}, OUT_3_3);
	wire [3:0] OUT_3_4;
	CAS CAS_3_4( {OUT_3_3[0], OUT_2_3[1], M[4], Q[29]}, OUT_3_4);
	wire [3:0] OUT_3_5;
	CAS CAS_3_5( {OUT_3_4[0], OUT_2_4[1], M[5], Q[29]}, OUT_3_5);
	wire [3:0] OUT_3_6;
	CAS CAS_3_6( {OUT_3_5[0], OUT_2_5[1], M[6], Q[29]}, OUT_3_6);
	wire [3:0] OUT_3_7;
	CAS CAS_3_7( {OUT_3_6[0], OUT_2_6[1], M[7], Q[29]}, OUT_3_7);
	wire [3:0] OUT_3_8;
	CAS CAS_3_8( {OUT_3_7[0], OUT_2_7[1], M[8], Q[29]}, OUT_3_8);
	wire [3:0] OUT_3_9;
	CAS CAS_3_9( {OUT_3_8[0], OUT_2_8[1], M[9], Q[29]}, OUT_3_9);
	wire [3:0] OUT_3_10;
	CAS CAS_3_10( {OUT_3_9[0], OUT_2_9[1], M[10], Q[29]}, OUT_3_10);
	wire [3:0] OUT_3_11;
	CAS CAS_3_11( {OUT_3_10[0], OUT_2_10[1], M[11], Q[29]}, OUT_3_11);
	wire [3:0] OUT_3_12;
	CAS CAS_3_12( {OUT_3_11[0], OUT_2_11[1], M[12], Q[29]}, OUT_3_12);
	wire [3:0] OUT_3_13;
	CAS CAS_3_13( {OUT_3_12[0], OUT_2_12[1], M[13], Q[29]}, OUT_3_13);
	wire [3:0] OUT_3_14;
	CAS CAS_3_14( {OUT_3_13[0], OUT_2_13[1], M[14], Q[29]}, OUT_3_14);
	wire [3:0] OUT_3_15;
	CAS CAS_3_15( {OUT_3_14[0], OUT_2_14[1], M[15], Q[29]}, OUT_3_15);
	wire [3:0] OUT_3_16;
	CAS CAS_3_16( {OUT_3_15[0], OUT_2_15[1], M[16], Q[29]}, OUT_3_16);
	wire [3:0] OUT_3_17;
	CAS CAS_3_17( {OUT_3_16[0], OUT_2_16[1], M[17], Q[29]}, OUT_3_17);
	wire [3:0] OUT_3_18;
	CAS CAS_3_18( {OUT_3_17[0], OUT_2_17[1], M[18], Q[29]}, OUT_3_18);
	wire [3:0] OUT_3_19;
	CAS CAS_3_19( {OUT_3_18[0], OUT_2_18[1], M[19], Q[29]}, OUT_3_19);
	wire [3:0] OUT_3_20;
	CAS CAS_3_20( {OUT_3_19[0], OUT_2_19[1], M[20], Q[29]}, OUT_3_20);
	wire [3:0] OUT_3_21;
	CAS CAS_3_21( {OUT_3_20[0], OUT_2_20[1], M[21], Q[29]}, OUT_3_21);
	wire [3:0] OUT_3_22;
	CAS CAS_3_22( {OUT_3_21[0], OUT_2_21[1], M[22], Q[29]}, OUT_3_22);
	wire [3:0] OUT_3_23;
	CAS CAS_3_23( {OUT_3_22[0], OUT_2_22[1], M[23], Q[29]}, OUT_3_23);
	wire [3:0] OUT_3_24;
	CAS CAS_3_24( {OUT_3_23[0], OUT_2_23[1], M[24], Q[29]}, OUT_3_24);
	wire [3:0] OUT_3_25;
	CAS CAS_3_25( {OUT_3_24[0], OUT_2_24[1], M[25], Q[29]}, OUT_3_25);
	wire [3:0] OUT_3_26;
	CAS CAS_3_26( {OUT_3_25[0], OUT_2_25[1], M[26], Q[29]}, OUT_3_26);
	wire [3:0] OUT_3_27;
	CAS CAS_3_27( {OUT_3_26[0], OUT_2_26[1], M[27], Q[29]}, OUT_3_27);
	wire [3:0] OUT_3_28;
	CAS CAS_3_28( {OUT_3_27[0], OUT_2_27[1], M[28], Q[29]}, OUT_3_28);
	wire [3:0] OUT_3_29;
	CAS CAS_3_29( {OUT_3_28[0], OUT_2_28[1], M[29], Q[29]}, OUT_3_29);
	wire [3:0] OUT_3_30;
	CAS CAS_3_30( {OUT_3_29[0], OUT_2_29[1], M[30], Q[29]}, OUT_3_30);
	wire [3:0] OUT_3_31;
	CAS CAS_3_31( {OUT_3_30[0], OUT_2_30[1], M[31], Q[29]}, OUT_3_31);
	assign Q[28] = OUT_3_31[0];

// Level - 5
	wire [3:0] OUT_4_0;
	CAS CAS_4_0( {Q[28], D[27], M[0], Q[28]}, OUT_4_0);
	wire [3:0] OUT_4_1;
	CAS CAS_4_1( {OUT_4_0[0], OUT_3_0[1], M[1], Q[28]}, OUT_4_1);
	wire [3:0] OUT_4_2;
	CAS CAS_4_2( {OUT_4_1[0], OUT_3_1[1], M[2], Q[28]}, OUT_4_2);
	wire [3:0] OUT_4_3;
	CAS CAS_4_3( {OUT_4_2[0], OUT_3_2[1], M[3], Q[28]}, OUT_4_3);
	wire [3:0] OUT_4_4;
	CAS CAS_4_4( {OUT_4_3[0], OUT_3_3[1], M[4], Q[28]}, OUT_4_4);
	wire [3:0] OUT_4_5;
	CAS CAS_4_5( {OUT_4_4[0], OUT_3_4[1], M[5], Q[28]}, OUT_4_5);
	wire [3:0] OUT_4_6;
	CAS CAS_4_6( {OUT_4_5[0], OUT_3_5[1], M[6], Q[28]}, OUT_4_6);
	wire [3:0] OUT_4_7;
	CAS CAS_4_7( {OUT_4_6[0], OUT_3_6[1], M[7], Q[28]}, OUT_4_7);
	wire [3:0] OUT_4_8;
	CAS CAS_4_8( {OUT_4_7[0], OUT_3_7[1], M[8], Q[28]}, OUT_4_8);
	wire [3:0] OUT_4_9;
	CAS CAS_4_9( {OUT_4_8[0], OUT_3_8[1], M[9], Q[28]}, OUT_4_9);
	wire [3:0] OUT_4_10;
	CAS CAS_4_10( {OUT_4_9[0], OUT_3_9[1], M[10], Q[28]}, OUT_4_10);
	wire [3:0] OUT_4_11;
	CAS CAS_4_11( {OUT_4_10[0], OUT_3_10[1], M[11], Q[28]}, OUT_4_11);
	wire [3:0] OUT_4_12;
	CAS CAS_4_12( {OUT_4_11[0], OUT_3_11[1], M[12], Q[28]}, OUT_4_12);
	wire [3:0] OUT_4_13;
	CAS CAS_4_13( {OUT_4_12[0], OUT_3_12[1], M[13], Q[28]}, OUT_4_13);
	wire [3:0] OUT_4_14;
	CAS CAS_4_14( {OUT_4_13[0], OUT_3_13[1], M[14], Q[28]}, OUT_4_14);
	wire [3:0] OUT_4_15;
	CAS CAS_4_15( {OUT_4_14[0], OUT_3_14[1], M[15], Q[28]}, OUT_4_15);
	wire [3:0] OUT_4_16;
	CAS CAS_4_16( {OUT_4_15[0], OUT_3_15[1], M[16], Q[28]}, OUT_4_16);
	wire [3:0] OUT_4_17;
	CAS CAS_4_17( {OUT_4_16[0], OUT_3_16[1], M[17], Q[28]}, OUT_4_17);
	wire [3:0] OUT_4_18;
	CAS CAS_4_18( {OUT_4_17[0], OUT_3_17[1], M[18], Q[28]}, OUT_4_18);
	wire [3:0] OUT_4_19;
	CAS CAS_4_19( {OUT_4_18[0], OUT_3_18[1], M[19], Q[28]}, OUT_4_19);
	wire [3:0] OUT_4_20;
	CAS CAS_4_20( {OUT_4_19[0], OUT_3_19[1], M[20], Q[28]}, OUT_4_20);
	wire [3:0] OUT_4_21;
	CAS CAS_4_21( {OUT_4_20[0], OUT_3_20[1], M[21], Q[28]}, OUT_4_21);
	wire [3:0] OUT_4_22;
	CAS CAS_4_22( {OUT_4_21[0], OUT_3_21[1], M[22], Q[28]}, OUT_4_22);
	wire [3:0] OUT_4_23;
	CAS CAS_4_23( {OUT_4_22[0], OUT_3_22[1], M[23], Q[28]}, OUT_4_23);
	wire [3:0] OUT_4_24;
	CAS CAS_4_24( {OUT_4_23[0], OUT_3_23[1], M[24], Q[28]}, OUT_4_24);
	wire [3:0] OUT_4_25;
	CAS CAS_4_25( {OUT_4_24[0], OUT_3_24[1], M[25], Q[28]}, OUT_4_25);
	wire [3:0] OUT_4_26;
	CAS CAS_4_26( {OUT_4_25[0], OUT_3_25[1], M[26], Q[28]}, OUT_4_26);
	wire [3:0] OUT_4_27;
	CAS CAS_4_27( {OUT_4_26[0], OUT_3_26[1], M[27], Q[28]}, OUT_4_27);
	wire [3:0] OUT_4_28;
	CAS CAS_4_28( {OUT_4_27[0], OUT_3_27[1], M[28], Q[28]}, OUT_4_28);
	wire [3:0] OUT_4_29;
	CAS CAS_4_29( {OUT_4_28[0], OUT_3_28[1], M[29], Q[28]}, OUT_4_29);
	wire [3:0] OUT_4_30;
	CAS CAS_4_30( {OUT_4_29[0], OUT_3_29[1], M[30], Q[28]}, OUT_4_30);
	wire [3:0] OUT_4_31;
	CAS CAS_4_31( {OUT_4_30[0], OUT_3_30[1], M[31], Q[28]}, OUT_4_31);
	assign Q[27] = OUT_4_31[0];

// Level - 6
	wire [3:0] OUT_5_0;
	CAS CAS_5_0( {Q[27], D[26], M[0], Q[27]}, OUT_5_0);
	wire [3:0] OUT_5_1;
	CAS CAS_5_1( {OUT_5_0[0], OUT_4_0[1], M[1], Q[27]}, OUT_5_1);
	wire [3:0] OUT_5_2;
	CAS CAS_5_2( {OUT_5_1[0], OUT_4_1[1], M[2], Q[27]}, OUT_5_2);
	wire [3:0] OUT_5_3;
	CAS CAS_5_3( {OUT_5_2[0], OUT_4_2[1], M[3], Q[27]}, OUT_5_3);
	wire [3:0] OUT_5_4;
	CAS CAS_5_4( {OUT_5_3[0], OUT_4_3[1], M[4], Q[27]}, OUT_5_4);
	wire [3:0] OUT_5_5;
	CAS CAS_5_5( {OUT_5_4[0], OUT_4_4[1], M[5], Q[27]}, OUT_5_5);
	wire [3:0] OUT_5_6;
	CAS CAS_5_6( {OUT_5_5[0], OUT_4_5[1], M[6], Q[27]}, OUT_5_6);
	wire [3:0] OUT_5_7;
	CAS CAS_5_7( {OUT_5_6[0], OUT_4_6[1], M[7], Q[27]}, OUT_5_7);
	wire [3:0] OUT_5_8;
	CAS CAS_5_8( {OUT_5_7[0], OUT_4_7[1], M[8], Q[27]}, OUT_5_8);
	wire [3:0] OUT_5_9;
	CAS CAS_5_9( {OUT_5_8[0], OUT_4_8[1], M[9], Q[27]}, OUT_5_9);
	wire [3:0] OUT_5_10;
	CAS CAS_5_10( {OUT_5_9[0], OUT_4_9[1], M[10], Q[27]}, OUT_5_10);
	wire [3:0] OUT_5_11;
	CAS CAS_5_11( {OUT_5_10[0], OUT_4_10[1], M[11], Q[27]}, OUT_5_11);
	wire [3:0] OUT_5_12;
	CAS CAS_5_12( {OUT_5_11[0], OUT_4_11[1], M[12], Q[27]}, OUT_5_12);
	wire [3:0] OUT_5_13;
	CAS CAS_5_13( {OUT_5_12[0], OUT_4_12[1], M[13], Q[27]}, OUT_5_13);
	wire [3:0] OUT_5_14;
	CAS CAS_5_14( {OUT_5_13[0], OUT_4_13[1], M[14], Q[27]}, OUT_5_14);
	wire [3:0] OUT_5_15;
	CAS CAS_5_15( {OUT_5_14[0], OUT_4_14[1], M[15], Q[27]}, OUT_5_15);
	wire [3:0] OUT_5_16;
	CAS CAS_5_16( {OUT_5_15[0], OUT_4_15[1], M[16], Q[27]}, OUT_5_16);
	wire [3:0] OUT_5_17;
	CAS CAS_5_17( {OUT_5_16[0], OUT_4_16[1], M[17], Q[27]}, OUT_5_17);
	wire [3:0] OUT_5_18;
	CAS CAS_5_18( {OUT_5_17[0], OUT_4_17[1], M[18], Q[27]}, OUT_5_18);
	wire [3:0] OUT_5_19;
	CAS CAS_5_19( {OUT_5_18[0], OUT_4_18[1], M[19], Q[27]}, OUT_5_19);
	wire [3:0] OUT_5_20;
	CAS CAS_5_20( {OUT_5_19[0], OUT_4_19[1], M[20], Q[27]}, OUT_5_20);
	wire [3:0] OUT_5_21;
	CAS CAS_5_21( {OUT_5_20[0], OUT_4_20[1], M[21], Q[27]}, OUT_5_21);
	wire [3:0] OUT_5_22;
	CAS CAS_5_22( {OUT_5_21[0], OUT_4_21[1], M[22], Q[27]}, OUT_5_22);
	wire [3:0] OUT_5_23;
	CAS CAS_5_23( {OUT_5_22[0], OUT_4_22[1], M[23], Q[27]}, OUT_5_23);
	wire [3:0] OUT_5_24;
	CAS CAS_5_24( {OUT_5_23[0], OUT_4_23[1], M[24], Q[27]}, OUT_5_24);
	wire [3:0] OUT_5_25;
	CAS CAS_5_25( {OUT_5_24[0], OUT_4_24[1], M[25], Q[27]}, OUT_5_25);
	wire [3:0] OUT_5_26;
	CAS CAS_5_26( {OUT_5_25[0], OUT_4_25[1], M[26], Q[27]}, OUT_5_26);
	wire [3:0] OUT_5_27;
	CAS CAS_5_27( {OUT_5_26[0], OUT_4_26[1], M[27], Q[27]}, OUT_5_27);
	wire [3:0] OUT_5_28;
	CAS CAS_5_28( {OUT_5_27[0], OUT_4_27[1], M[28], Q[27]}, OUT_5_28);
	wire [3:0] OUT_5_29;
	CAS CAS_5_29( {OUT_5_28[0], OUT_4_28[1], M[29], Q[27]}, OUT_5_29);
	wire [3:0] OUT_5_30;
	CAS CAS_5_30( {OUT_5_29[0], OUT_4_29[1], M[30], Q[27]}, OUT_5_30);
	wire [3:0] OUT_5_31;
	CAS CAS_5_31( {OUT_5_30[0], OUT_4_30[1], M[31], Q[27]}, OUT_5_31);
	assign Q[26] = OUT_5_31[0];

// Level - 7
	wire [3:0] OUT_6_0;
	CAS CAS_6_0( {Q[26], D[25], M[0], Q[26]}, OUT_6_0);
	wire [3:0] OUT_6_1;
	CAS CAS_6_1( {OUT_6_0[0], OUT_5_0[1], M[1], Q[26]}, OUT_6_1);
	wire [3:0] OUT_6_2;
	CAS CAS_6_2( {OUT_6_1[0], OUT_5_1[1], M[2], Q[26]}, OUT_6_2);
	wire [3:0] OUT_6_3;
	CAS CAS_6_3( {OUT_6_2[0], OUT_5_2[1], M[3], Q[26]}, OUT_6_3);
	wire [3:0] OUT_6_4;
	CAS CAS_6_4( {OUT_6_3[0], OUT_5_3[1], M[4], Q[26]}, OUT_6_4);
	wire [3:0] OUT_6_5;
	CAS CAS_6_5( {OUT_6_4[0], OUT_5_4[1], M[5], Q[26]}, OUT_6_5);
	wire [3:0] OUT_6_6;
	CAS CAS_6_6( {OUT_6_5[0], OUT_5_5[1], M[6], Q[26]}, OUT_6_6);
	wire [3:0] OUT_6_7;
	CAS CAS_6_7( {OUT_6_6[0], OUT_5_6[1], M[7], Q[26]}, OUT_6_7);
	wire [3:0] OUT_6_8;
	CAS CAS_6_8( {OUT_6_7[0], OUT_5_7[1], M[8], Q[26]}, OUT_6_8);
	wire [3:0] OUT_6_9;
	CAS CAS_6_9( {OUT_6_8[0], OUT_5_8[1], M[9], Q[26]}, OUT_6_9);
	wire [3:0] OUT_6_10;
	CAS CAS_6_10( {OUT_6_9[0], OUT_5_9[1], M[10], Q[26]}, OUT_6_10);
	wire [3:0] OUT_6_11;
	CAS CAS_6_11( {OUT_6_10[0], OUT_5_10[1], M[11], Q[26]}, OUT_6_11);
	wire [3:0] OUT_6_12;
	CAS CAS_6_12( {OUT_6_11[0], OUT_5_11[1], M[12], Q[26]}, OUT_6_12);
	wire [3:0] OUT_6_13;
	CAS CAS_6_13( {OUT_6_12[0], OUT_5_12[1], M[13], Q[26]}, OUT_6_13);
	wire [3:0] OUT_6_14;
	CAS CAS_6_14( {OUT_6_13[0], OUT_5_13[1], M[14], Q[26]}, OUT_6_14);
	wire [3:0] OUT_6_15;
	CAS CAS_6_15( {OUT_6_14[0], OUT_5_14[1], M[15], Q[26]}, OUT_6_15);
	wire [3:0] OUT_6_16;
	CAS CAS_6_16( {OUT_6_15[0], OUT_5_15[1], M[16], Q[26]}, OUT_6_16);
	wire [3:0] OUT_6_17;
	CAS CAS_6_17( {OUT_6_16[0], OUT_5_16[1], M[17], Q[26]}, OUT_6_17);
	wire [3:0] OUT_6_18;
	CAS CAS_6_18( {OUT_6_17[0], OUT_5_17[1], M[18], Q[26]}, OUT_6_18);
	wire [3:0] OUT_6_19;
	CAS CAS_6_19( {OUT_6_18[0], OUT_5_18[1], M[19], Q[26]}, OUT_6_19);
	wire [3:0] OUT_6_20;
	CAS CAS_6_20( {OUT_6_19[0], OUT_5_19[1], M[20], Q[26]}, OUT_6_20);
	wire [3:0] OUT_6_21;
	CAS CAS_6_21( {OUT_6_20[0], OUT_5_20[1], M[21], Q[26]}, OUT_6_21);
	wire [3:0] OUT_6_22;
	CAS CAS_6_22( {OUT_6_21[0], OUT_5_21[1], M[22], Q[26]}, OUT_6_22);
	wire [3:0] OUT_6_23;
	CAS CAS_6_23( {OUT_6_22[0], OUT_5_22[1], M[23], Q[26]}, OUT_6_23);
	wire [3:0] OUT_6_24;
	CAS CAS_6_24( {OUT_6_23[0], OUT_5_23[1], M[24], Q[26]}, OUT_6_24);
	wire [3:0] OUT_6_25;
	CAS CAS_6_25( {OUT_6_24[0], OUT_5_24[1], M[25], Q[26]}, OUT_6_25);
	wire [3:0] OUT_6_26;
	CAS CAS_6_26( {OUT_6_25[0], OUT_5_25[1], M[26], Q[26]}, OUT_6_26);
	wire [3:0] OUT_6_27;
	CAS CAS_6_27( {OUT_6_26[0], OUT_5_26[1], M[27], Q[26]}, OUT_6_27);
	wire [3:0] OUT_6_28;
	CAS CAS_6_28( {OUT_6_27[0], OUT_5_27[1], M[28], Q[26]}, OUT_6_28);
	wire [3:0] OUT_6_29;
	CAS CAS_6_29( {OUT_6_28[0], OUT_5_28[1], M[29], Q[26]}, OUT_6_29);
	wire [3:0] OUT_6_30;
	CAS CAS_6_30( {OUT_6_29[0], OUT_5_29[1], M[30], Q[26]}, OUT_6_30);
	wire [3:0] OUT_6_31;
	CAS CAS_6_31( {OUT_6_30[0], OUT_5_30[1], M[31], Q[26]}, OUT_6_31);
	assign Q[25] = OUT_6_31[0];

// Level - 8
	wire [3:0] OUT_7_0;
	CAS CAS_7_0( {Q[25], D[24], M[0], Q[25]}, OUT_7_0);
	wire [3:0] OUT_7_1;
	CAS CAS_7_1( {OUT_7_0[0], OUT_6_0[1], M[1], Q[25]}, OUT_7_1);
	wire [3:0] OUT_7_2;
	CAS CAS_7_2( {OUT_7_1[0], OUT_6_1[1], M[2], Q[25]}, OUT_7_2);
	wire [3:0] OUT_7_3;
	CAS CAS_7_3( {OUT_7_2[0], OUT_6_2[1], M[3], Q[25]}, OUT_7_3);
	wire [3:0] OUT_7_4;
	CAS CAS_7_4( {OUT_7_3[0], OUT_6_3[1], M[4], Q[25]}, OUT_7_4);
	wire [3:0] OUT_7_5;
	CAS CAS_7_5( {OUT_7_4[0], OUT_6_4[1], M[5], Q[25]}, OUT_7_5);
	wire [3:0] OUT_7_6;
	CAS CAS_7_6( {OUT_7_5[0], OUT_6_5[1], M[6], Q[25]}, OUT_7_6);
	wire [3:0] OUT_7_7;
	CAS CAS_7_7( {OUT_7_6[0], OUT_6_6[1], M[7], Q[25]}, OUT_7_7);
	wire [3:0] OUT_7_8;
	CAS CAS_7_8( {OUT_7_7[0], OUT_6_7[1], M[8], Q[25]}, OUT_7_8);
	wire [3:0] OUT_7_9;
	CAS CAS_7_9( {OUT_7_8[0], OUT_6_8[1], M[9], Q[25]}, OUT_7_9);
	wire [3:0] OUT_7_10;
	CAS CAS_7_10( {OUT_7_9[0], OUT_6_9[1], M[10], Q[25]}, OUT_7_10);
	wire [3:0] OUT_7_11;
	CAS CAS_7_11( {OUT_7_10[0], OUT_6_10[1], M[11], Q[25]}, OUT_7_11);
	wire [3:0] OUT_7_12;
	CAS CAS_7_12( {OUT_7_11[0], OUT_6_11[1], M[12], Q[25]}, OUT_7_12);
	wire [3:0] OUT_7_13;
	CAS CAS_7_13( {OUT_7_12[0], OUT_6_12[1], M[13], Q[25]}, OUT_7_13);
	wire [3:0] OUT_7_14;
	CAS CAS_7_14( {OUT_7_13[0], OUT_6_13[1], M[14], Q[25]}, OUT_7_14);
	wire [3:0] OUT_7_15;
	CAS CAS_7_15( {OUT_7_14[0], OUT_6_14[1], M[15], Q[25]}, OUT_7_15);
	wire [3:0] OUT_7_16;
	CAS CAS_7_16( {OUT_7_15[0], OUT_6_15[1], M[16], Q[25]}, OUT_7_16);
	wire [3:0] OUT_7_17;
	CAS CAS_7_17( {OUT_7_16[0], OUT_6_16[1], M[17], Q[25]}, OUT_7_17);
	wire [3:0] OUT_7_18;
	CAS CAS_7_18( {OUT_7_17[0], OUT_6_17[1], M[18], Q[25]}, OUT_7_18);
	wire [3:0] OUT_7_19;
	CAS CAS_7_19( {OUT_7_18[0], OUT_6_18[1], M[19], Q[25]}, OUT_7_19);
	wire [3:0] OUT_7_20;
	CAS CAS_7_20( {OUT_7_19[0], OUT_6_19[1], M[20], Q[25]}, OUT_7_20);
	wire [3:0] OUT_7_21;
	CAS CAS_7_21( {OUT_7_20[0], OUT_6_20[1], M[21], Q[25]}, OUT_7_21);
	wire [3:0] OUT_7_22;
	CAS CAS_7_22( {OUT_7_21[0], OUT_6_21[1], M[22], Q[25]}, OUT_7_22);
	wire [3:0] OUT_7_23;
	CAS CAS_7_23( {OUT_7_22[0], OUT_6_22[1], M[23], Q[25]}, OUT_7_23);
	wire [3:0] OUT_7_24;
	CAS CAS_7_24( {OUT_7_23[0], OUT_6_23[1], M[24], Q[25]}, OUT_7_24);
	wire [3:0] OUT_7_25;
	CAS CAS_7_25( {OUT_7_24[0], OUT_6_24[1], M[25], Q[25]}, OUT_7_25);
	wire [3:0] OUT_7_26;
	CAS CAS_7_26( {OUT_7_25[0], OUT_6_25[1], M[26], Q[25]}, OUT_7_26);
	wire [3:0] OUT_7_27;
	CAS CAS_7_27( {OUT_7_26[0], OUT_6_26[1], M[27], Q[25]}, OUT_7_27);
	wire [3:0] OUT_7_28;
	CAS CAS_7_28( {OUT_7_27[0], OUT_6_27[1], M[28], Q[25]}, OUT_7_28);
	wire [3:0] OUT_7_29;
	CAS CAS_7_29( {OUT_7_28[0], OUT_6_28[1], M[29], Q[25]}, OUT_7_29);
	wire [3:0] OUT_7_30;
	CAS CAS_7_30( {OUT_7_29[0], OUT_6_29[1], M[30], Q[25]}, OUT_7_30);
	wire [3:0] OUT_7_31;
	CAS CAS_7_31( {OUT_7_30[0], OUT_6_30[1], M[31], Q[25]}, OUT_7_31);
	assign Q[24] = OUT_7_31[0];

// Level - 9
	wire [3:0] OUT_8_0;
	CAS CAS_8_0( {Q[24], D[23], M[0], Q[24]}, OUT_8_0);
	wire [3:0] OUT_8_1;
	CAS CAS_8_1( {OUT_8_0[0], OUT_7_0[1], M[1], Q[24]}, OUT_8_1);
	wire [3:0] OUT_8_2;
	CAS CAS_8_2( {OUT_8_1[0], OUT_7_1[1], M[2], Q[24]}, OUT_8_2);
	wire [3:0] OUT_8_3;
	CAS CAS_8_3( {OUT_8_2[0], OUT_7_2[1], M[3], Q[24]}, OUT_8_3);
	wire [3:0] OUT_8_4;
	CAS CAS_8_4( {OUT_8_3[0], OUT_7_3[1], M[4], Q[24]}, OUT_8_4);
	wire [3:0] OUT_8_5;
	CAS CAS_8_5( {OUT_8_4[0], OUT_7_4[1], M[5], Q[24]}, OUT_8_5);
	wire [3:0] OUT_8_6;
	CAS CAS_8_6( {OUT_8_5[0], OUT_7_5[1], M[6], Q[24]}, OUT_8_6);
	wire [3:0] OUT_8_7;
	CAS CAS_8_7( {OUT_8_6[0], OUT_7_6[1], M[7], Q[24]}, OUT_8_7);
	wire [3:0] OUT_8_8;
	CAS CAS_8_8( {OUT_8_7[0], OUT_7_7[1], M[8], Q[24]}, OUT_8_8);
	wire [3:0] OUT_8_9;
	CAS CAS_8_9( {OUT_8_8[0], OUT_7_8[1], M[9], Q[24]}, OUT_8_9);
	wire [3:0] OUT_8_10;
	CAS CAS_8_10( {OUT_8_9[0], OUT_7_9[1], M[10], Q[24]}, OUT_8_10);
	wire [3:0] OUT_8_11;
	CAS CAS_8_11( {OUT_8_10[0], OUT_7_10[1], M[11], Q[24]}, OUT_8_11);
	wire [3:0] OUT_8_12;
	CAS CAS_8_12( {OUT_8_11[0], OUT_7_11[1], M[12], Q[24]}, OUT_8_12);
	wire [3:0] OUT_8_13;
	CAS CAS_8_13( {OUT_8_12[0], OUT_7_12[1], M[13], Q[24]}, OUT_8_13);
	wire [3:0] OUT_8_14;
	CAS CAS_8_14( {OUT_8_13[0], OUT_7_13[1], M[14], Q[24]}, OUT_8_14);
	wire [3:0] OUT_8_15;
	CAS CAS_8_15( {OUT_8_14[0], OUT_7_14[1], M[15], Q[24]}, OUT_8_15);
	wire [3:0] OUT_8_16;
	CAS CAS_8_16( {OUT_8_15[0], OUT_7_15[1], M[16], Q[24]}, OUT_8_16);
	wire [3:0] OUT_8_17;
	CAS CAS_8_17( {OUT_8_16[0], OUT_7_16[1], M[17], Q[24]}, OUT_8_17);
	wire [3:0] OUT_8_18;
	CAS CAS_8_18( {OUT_8_17[0], OUT_7_17[1], M[18], Q[24]}, OUT_8_18);
	wire [3:0] OUT_8_19;
	CAS CAS_8_19( {OUT_8_18[0], OUT_7_18[1], M[19], Q[24]}, OUT_8_19);
	wire [3:0] OUT_8_20;
	CAS CAS_8_20( {OUT_8_19[0], OUT_7_19[1], M[20], Q[24]}, OUT_8_20);
	wire [3:0] OUT_8_21;
	CAS CAS_8_21( {OUT_8_20[0], OUT_7_20[1], M[21], Q[24]}, OUT_8_21);
	wire [3:0] OUT_8_22;
	CAS CAS_8_22( {OUT_8_21[0], OUT_7_21[1], M[22], Q[24]}, OUT_8_22);
	wire [3:0] OUT_8_23;
	CAS CAS_8_23( {OUT_8_22[0], OUT_7_22[1], M[23], Q[24]}, OUT_8_23);
	wire [3:0] OUT_8_24;
	CAS CAS_8_24( {OUT_8_23[0], OUT_7_23[1], M[24], Q[24]}, OUT_8_24);
	wire [3:0] OUT_8_25;
	CAS CAS_8_25( {OUT_8_24[0], OUT_7_24[1], M[25], Q[24]}, OUT_8_25);
	wire [3:0] OUT_8_26;
	CAS CAS_8_26( {OUT_8_25[0], OUT_7_25[1], M[26], Q[24]}, OUT_8_26);
	wire [3:0] OUT_8_27;
	CAS CAS_8_27( {OUT_8_26[0], OUT_7_26[1], M[27], Q[24]}, OUT_8_27);
	wire [3:0] OUT_8_28;
	CAS CAS_8_28( {OUT_8_27[0], OUT_7_27[1], M[28], Q[24]}, OUT_8_28);
	wire [3:0] OUT_8_29;
	CAS CAS_8_29( {OUT_8_28[0], OUT_7_28[1], M[29], Q[24]}, OUT_8_29);
	wire [3:0] OUT_8_30;
	CAS CAS_8_30( {OUT_8_29[0], OUT_7_29[1], M[30], Q[24]}, OUT_8_30);
	wire [3:0] OUT_8_31;
	CAS CAS_8_31( {OUT_8_30[0], OUT_7_30[1], M[31], Q[24]}, OUT_8_31);
	assign Q[23] = OUT_8_31[0];

// Level - 10
	wire [3:0] OUT_9_0;
	CAS CAS_9_0( {Q[23], D[22], M[0], Q[23]}, OUT_9_0);
	wire [3:0] OUT_9_1;
	CAS CAS_9_1( {OUT_9_0[0], OUT_8_0[1], M[1], Q[23]}, OUT_9_1);
	wire [3:0] OUT_9_2;
	CAS CAS_9_2( {OUT_9_1[0], OUT_8_1[1], M[2], Q[23]}, OUT_9_2);
	wire [3:0] OUT_9_3;
	CAS CAS_9_3( {OUT_9_2[0], OUT_8_2[1], M[3], Q[23]}, OUT_9_3);
	wire [3:0] OUT_9_4;
	CAS CAS_9_4( {OUT_9_3[0], OUT_8_3[1], M[4], Q[23]}, OUT_9_4);
	wire [3:0] OUT_9_5;
	CAS CAS_9_5( {OUT_9_4[0], OUT_8_4[1], M[5], Q[23]}, OUT_9_5);
	wire [3:0] OUT_9_6;
	CAS CAS_9_6( {OUT_9_5[0], OUT_8_5[1], M[6], Q[23]}, OUT_9_6);
	wire [3:0] OUT_9_7;
	CAS CAS_9_7( {OUT_9_6[0], OUT_8_6[1], M[7], Q[23]}, OUT_9_7);
	wire [3:0] OUT_9_8;
	CAS CAS_9_8( {OUT_9_7[0], OUT_8_7[1], M[8], Q[23]}, OUT_9_8);
	wire [3:0] OUT_9_9;
	CAS CAS_9_9( {OUT_9_8[0], OUT_8_8[1], M[9], Q[23]}, OUT_9_9);
	wire [3:0] OUT_9_10;
	CAS CAS_9_10( {OUT_9_9[0], OUT_8_9[1], M[10], Q[23]}, OUT_9_10);
	wire [3:0] OUT_9_11;
	CAS CAS_9_11( {OUT_9_10[0], OUT_8_10[1], M[11], Q[23]}, OUT_9_11);
	wire [3:0] OUT_9_12;
	CAS CAS_9_12( {OUT_9_11[0], OUT_8_11[1], M[12], Q[23]}, OUT_9_12);
	wire [3:0] OUT_9_13;
	CAS CAS_9_13( {OUT_9_12[0], OUT_8_12[1], M[13], Q[23]}, OUT_9_13);
	wire [3:0] OUT_9_14;
	CAS CAS_9_14( {OUT_9_13[0], OUT_8_13[1], M[14], Q[23]}, OUT_9_14);
	wire [3:0] OUT_9_15;
	CAS CAS_9_15( {OUT_9_14[0], OUT_8_14[1], M[15], Q[23]}, OUT_9_15);
	wire [3:0] OUT_9_16;
	CAS CAS_9_16( {OUT_9_15[0], OUT_8_15[1], M[16], Q[23]}, OUT_9_16);
	wire [3:0] OUT_9_17;
	CAS CAS_9_17( {OUT_9_16[0], OUT_8_16[1], M[17], Q[23]}, OUT_9_17);
	wire [3:0] OUT_9_18;
	CAS CAS_9_18( {OUT_9_17[0], OUT_8_17[1], M[18], Q[23]}, OUT_9_18);
	wire [3:0] OUT_9_19;
	CAS CAS_9_19( {OUT_9_18[0], OUT_8_18[1], M[19], Q[23]}, OUT_9_19);
	wire [3:0] OUT_9_20;
	CAS CAS_9_20( {OUT_9_19[0], OUT_8_19[1], M[20], Q[23]}, OUT_9_20);
	wire [3:0] OUT_9_21;
	CAS CAS_9_21( {OUT_9_20[0], OUT_8_20[1], M[21], Q[23]}, OUT_9_21);
	wire [3:0] OUT_9_22;
	CAS CAS_9_22( {OUT_9_21[0], OUT_8_21[1], M[22], Q[23]}, OUT_9_22);
	wire [3:0] OUT_9_23;
	CAS CAS_9_23( {OUT_9_22[0], OUT_8_22[1], M[23], Q[23]}, OUT_9_23);
	wire [3:0] OUT_9_24;
	CAS CAS_9_24( {OUT_9_23[0], OUT_8_23[1], M[24], Q[23]}, OUT_9_24);
	wire [3:0] OUT_9_25;
	CAS CAS_9_25( {OUT_9_24[0], OUT_8_24[1], M[25], Q[23]}, OUT_9_25);
	wire [3:0] OUT_9_26;
	CAS CAS_9_26( {OUT_9_25[0], OUT_8_25[1], M[26], Q[23]}, OUT_9_26);
	wire [3:0] OUT_9_27;
	CAS CAS_9_27( {OUT_9_26[0], OUT_8_26[1], M[27], Q[23]}, OUT_9_27);
	wire [3:0] OUT_9_28;
	CAS CAS_9_28( {OUT_9_27[0], OUT_8_27[1], M[28], Q[23]}, OUT_9_28);
	wire [3:0] OUT_9_29;
	CAS CAS_9_29( {OUT_9_28[0], OUT_8_28[1], M[29], Q[23]}, OUT_9_29);
	wire [3:0] OUT_9_30;
	CAS CAS_9_30( {OUT_9_29[0], OUT_8_29[1], M[30], Q[23]}, OUT_9_30);
	wire [3:0] OUT_9_31;
	CAS CAS_9_31( {OUT_9_30[0], OUT_8_30[1], M[31], Q[23]}, OUT_9_31);
	assign Q[22] = OUT_9_31[0];

// Level - 11
	wire [3:0] OUT_10_0;
	CAS CAS_10_0( {Q[22], D[21], M[0], Q[22]}, OUT_10_0);
	wire [3:0] OUT_10_1;
	CAS CAS_10_1( {OUT_10_0[0], OUT_9_0[1], M[1], Q[22]}, OUT_10_1);
	wire [3:0] OUT_10_2;
	CAS CAS_10_2( {OUT_10_1[0], OUT_9_1[1], M[2], Q[22]}, OUT_10_2);
	wire [3:0] OUT_10_3;
	CAS CAS_10_3( {OUT_10_2[0], OUT_9_2[1], M[3], Q[22]}, OUT_10_3);
	wire [3:0] OUT_10_4;
	CAS CAS_10_4( {OUT_10_3[0], OUT_9_3[1], M[4], Q[22]}, OUT_10_4);
	wire [3:0] OUT_10_5;
	CAS CAS_10_5( {OUT_10_4[0], OUT_9_4[1], M[5], Q[22]}, OUT_10_5);
	wire [3:0] OUT_10_6;
	CAS CAS_10_6( {OUT_10_5[0], OUT_9_5[1], M[6], Q[22]}, OUT_10_6);
	wire [3:0] OUT_10_7;
	CAS CAS_10_7( {OUT_10_6[0], OUT_9_6[1], M[7], Q[22]}, OUT_10_7);
	wire [3:0] OUT_10_8;
	CAS CAS_10_8( {OUT_10_7[0], OUT_9_7[1], M[8], Q[22]}, OUT_10_8);
	wire [3:0] OUT_10_9;
	CAS CAS_10_9( {OUT_10_8[0], OUT_9_8[1], M[9], Q[22]}, OUT_10_9);
	wire [3:0] OUT_10_10;
	CAS CAS_10_10( {OUT_10_9[0], OUT_9_9[1], M[10], Q[22]}, OUT_10_10);
	wire [3:0] OUT_10_11;
	CAS CAS_10_11( {OUT_10_10[0], OUT_9_10[1], M[11], Q[22]}, OUT_10_11);
	wire [3:0] OUT_10_12;
	CAS CAS_10_12( {OUT_10_11[0], OUT_9_11[1], M[12], Q[22]}, OUT_10_12);
	wire [3:0] OUT_10_13;
	CAS CAS_10_13( {OUT_10_12[0], OUT_9_12[1], M[13], Q[22]}, OUT_10_13);
	wire [3:0] OUT_10_14;
	CAS CAS_10_14( {OUT_10_13[0], OUT_9_13[1], M[14], Q[22]}, OUT_10_14);
	wire [3:0] OUT_10_15;
	CAS CAS_10_15( {OUT_10_14[0], OUT_9_14[1], M[15], Q[22]}, OUT_10_15);
	wire [3:0] OUT_10_16;
	CAS CAS_10_16( {OUT_10_15[0], OUT_9_15[1], M[16], Q[22]}, OUT_10_16);
	wire [3:0] OUT_10_17;
	CAS CAS_10_17( {OUT_10_16[0], OUT_9_16[1], M[17], Q[22]}, OUT_10_17);
	wire [3:0] OUT_10_18;
	CAS CAS_10_18( {OUT_10_17[0], OUT_9_17[1], M[18], Q[22]}, OUT_10_18);
	wire [3:0] OUT_10_19;
	CAS CAS_10_19( {OUT_10_18[0], OUT_9_18[1], M[19], Q[22]}, OUT_10_19);
	wire [3:0] OUT_10_20;
	CAS CAS_10_20( {OUT_10_19[0], OUT_9_19[1], M[20], Q[22]}, OUT_10_20);
	wire [3:0] OUT_10_21;
	CAS CAS_10_21( {OUT_10_20[0], OUT_9_20[1], M[21], Q[22]}, OUT_10_21);
	wire [3:0] OUT_10_22;
	CAS CAS_10_22( {OUT_10_21[0], OUT_9_21[1], M[22], Q[22]}, OUT_10_22);
	wire [3:0] OUT_10_23;
	CAS CAS_10_23( {OUT_10_22[0], OUT_9_22[1], M[23], Q[22]}, OUT_10_23);
	wire [3:0] OUT_10_24;
	CAS CAS_10_24( {OUT_10_23[0], OUT_9_23[1], M[24], Q[22]}, OUT_10_24);
	wire [3:0] OUT_10_25;
	CAS CAS_10_25( {OUT_10_24[0], OUT_9_24[1], M[25], Q[22]}, OUT_10_25);
	wire [3:0] OUT_10_26;
	CAS CAS_10_26( {OUT_10_25[0], OUT_9_25[1], M[26], Q[22]}, OUT_10_26);
	wire [3:0] OUT_10_27;
	CAS CAS_10_27( {OUT_10_26[0], OUT_9_26[1], M[27], Q[22]}, OUT_10_27);
	wire [3:0] OUT_10_28;
	CAS CAS_10_28( {OUT_10_27[0], OUT_9_27[1], M[28], Q[22]}, OUT_10_28);
	wire [3:0] OUT_10_29;
	CAS CAS_10_29( {OUT_10_28[0], OUT_9_28[1], M[29], Q[22]}, OUT_10_29);
	wire [3:0] OUT_10_30;
	CAS CAS_10_30( {OUT_10_29[0], OUT_9_29[1], M[30], Q[22]}, OUT_10_30);
	wire [3:0] OUT_10_31;
	CAS CAS_10_31( {OUT_10_30[0], OUT_9_30[1], M[31], Q[22]}, OUT_10_31);
	assign Q[21] = OUT_10_31[0];

// Level - 12
	wire [3:0] OUT_11_0;
	CAS CAS_11_0( {Q[21], D[20], M[0], Q[21]}, OUT_11_0);
	wire [3:0] OUT_11_1;
	CAS CAS_11_1( {OUT_11_0[0], OUT_10_0[1], M[1], Q[21]}, OUT_11_1);
	wire [3:0] OUT_11_2;
	CAS CAS_11_2( {OUT_11_1[0], OUT_10_1[1], M[2], Q[21]}, OUT_11_2);
	wire [3:0] OUT_11_3;
	CAS CAS_11_3( {OUT_11_2[0], OUT_10_2[1], M[3], Q[21]}, OUT_11_3);
	wire [3:0] OUT_11_4;
	CAS CAS_11_4( {OUT_11_3[0], OUT_10_3[1], M[4], Q[21]}, OUT_11_4);
	wire [3:0] OUT_11_5;
	CAS CAS_11_5( {OUT_11_4[0], OUT_10_4[1], M[5], Q[21]}, OUT_11_5);
	wire [3:0] OUT_11_6;
	CAS CAS_11_6( {OUT_11_5[0], OUT_10_5[1], M[6], Q[21]}, OUT_11_6);
	wire [3:0] OUT_11_7;
	CAS CAS_11_7( {OUT_11_6[0], OUT_10_6[1], M[7], Q[21]}, OUT_11_7);
	wire [3:0] OUT_11_8;
	CAS CAS_11_8( {OUT_11_7[0], OUT_10_7[1], M[8], Q[21]}, OUT_11_8);
	wire [3:0] OUT_11_9;
	CAS CAS_11_9( {OUT_11_8[0], OUT_10_8[1], M[9], Q[21]}, OUT_11_9);
	wire [3:0] OUT_11_10;
	CAS CAS_11_10( {OUT_11_9[0], OUT_10_9[1], M[10], Q[21]}, OUT_11_10);
	wire [3:0] OUT_11_11;
	CAS CAS_11_11( {OUT_11_10[0], OUT_10_10[1], M[11], Q[21]}, OUT_11_11);
	wire [3:0] OUT_11_12;
	CAS CAS_11_12( {OUT_11_11[0], OUT_10_11[1], M[12], Q[21]}, OUT_11_12);
	wire [3:0] OUT_11_13;
	CAS CAS_11_13( {OUT_11_12[0], OUT_10_12[1], M[13], Q[21]}, OUT_11_13);
	wire [3:0] OUT_11_14;
	CAS CAS_11_14( {OUT_11_13[0], OUT_10_13[1], M[14], Q[21]}, OUT_11_14);
	wire [3:0] OUT_11_15;
	CAS CAS_11_15( {OUT_11_14[0], OUT_10_14[1], M[15], Q[21]}, OUT_11_15);
	wire [3:0] OUT_11_16;
	CAS CAS_11_16( {OUT_11_15[0], OUT_10_15[1], M[16], Q[21]}, OUT_11_16);
	wire [3:0] OUT_11_17;
	CAS CAS_11_17( {OUT_11_16[0], OUT_10_16[1], M[17], Q[21]}, OUT_11_17);
	wire [3:0] OUT_11_18;
	CAS CAS_11_18( {OUT_11_17[0], OUT_10_17[1], M[18], Q[21]}, OUT_11_18);
	wire [3:0] OUT_11_19;
	CAS CAS_11_19( {OUT_11_18[0], OUT_10_18[1], M[19], Q[21]}, OUT_11_19);
	wire [3:0] OUT_11_20;
	CAS CAS_11_20( {OUT_11_19[0], OUT_10_19[1], M[20], Q[21]}, OUT_11_20);
	wire [3:0] OUT_11_21;
	CAS CAS_11_21( {OUT_11_20[0], OUT_10_20[1], M[21], Q[21]}, OUT_11_21);
	wire [3:0] OUT_11_22;
	CAS CAS_11_22( {OUT_11_21[0], OUT_10_21[1], M[22], Q[21]}, OUT_11_22);
	wire [3:0] OUT_11_23;
	CAS CAS_11_23( {OUT_11_22[0], OUT_10_22[1], M[23], Q[21]}, OUT_11_23);
	wire [3:0] OUT_11_24;
	CAS CAS_11_24( {OUT_11_23[0], OUT_10_23[1], M[24], Q[21]}, OUT_11_24);
	wire [3:0] OUT_11_25;
	CAS CAS_11_25( {OUT_11_24[0], OUT_10_24[1], M[25], Q[21]}, OUT_11_25);
	wire [3:0] OUT_11_26;
	CAS CAS_11_26( {OUT_11_25[0], OUT_10_25[1], M[26], Q[21]}, OUT_11_26);
	wire [3:0] OUT_11_27;
	CAS CAS_11_27( {OUT_11_26[0], OUT_10_26[1], M[27], Q[21]}, OUT_11_27);
	wire [3:0] OUT_11_28;
	CAS CAS_11_28( {OUT_11_27[0], OUT_10_27[1], M[28], Q[21]}, OUT_11_28);
	wire [3:0] OUT_11_29;
	CAS CAS_11_29( {OUT_11_28[0], OUT_10_28[1], M[29], Q[21]}, OUT_11_29);
	wire [3:0] OUT_11_30;
	CAS CAS_11_30( {OUT_11_29[0], OUT_10_29[1], M[30], Q[21]}, OUT_11_30);
	wire [3:0] OUT_11_31;
	CAS CAS_11_31( {OUT_11_30[0], OUT_10_30[1], M[31], Q[21]}, OUT_11_31);
	assign Q[20] = OUT_11_31[0];

// Level - 13
	wire [3:0] OUT_12_0;
	CAS CAS_12_0( {Q[20], D[19], M[0], Q[20]}, OUT_12_0);
	wire [3:0] OUT_12_1;
	CAS CAS_12_1( {OUT_12_0[0], OUT_11_0[1], M[1], Q[20]}, OUT_12_1);
	wire [3:0] OUT_12_2;
	CAS CAS_12_2( {OUT_12_1[0], OUT_11_1[1], M[2], Q[20]}, OUT_12_2);
	wire [3:0] OUT_12_3;
	CAS CAS_12_3( {OUT_12_2[0], OUT_11_2[1], M[3], Q[20]}, OUT_12_3);
	wire [3:0] OUT_12_4;
	CAS CAS_12_4( {OUT_12_3[0], OUT_11_3[1], M[4], Q[20]}, OUT_12_4);
	wire [3:0] OUT_12_5;
	CAS CAS_12_5( {OUT_12_4[0], OUT_11_4[1], M[5], Q[20]}, OUT_12_5);
	wire [3:0] OUT_12_6;
	CAS CAS_12_6( {OUT_12_5[0], OUT_11_5[1], M[6], Q[20]}, OUT_12_6);
	wire [3:0] OUT_12_7;
	CAS CAS_12_7( {OUT_12_6[0], OUT_11_6[1], M[7], Q[20]}, OUT_12_7);
	wire [3:0] OUT_12_8;
	CAS CAS_12_8( {OUT_12_7[0], OUT_11_7[1], M[8], Q[20]}, OUT_12_8);
	wire [3:0] OUT_12_9;
	CAS CAS_12_9( {OUT_12_8[0], OUT_11_8[1], M[9], Q[20]}, OUT_12_9);
	wire [3:0] OUT_12_10;
	CAS CAS_12_10( {OUT_12_9[0], OUT_11_9[1], M[10], Q[20]}, OUT_12_10);
	wire [3:0] OUT_12_11;
	CAS CAS_12_11( {OUT_12_10[0], OUT_11_10[1], M[11], Q[20]}, OUT_12_11);
	wire [3:0] OUT_12_12;
	CAS CAS_12_12( {OUT_12_11[0], OUT_11_11[1], M[12], Q[20]}, OUT_12_12);
	wire [3:0] OUT_12_13;
	CAS CAS_12_13( {OUT_12_12[0], OUT_11_12[1], M[13], Q[20]}, OUT_12_13);
	wire [3:0] OUT_12_14;
	CAS CAS_12_14( {OUT_12_13[0], OUT_11_13[1], M[14], Q[20]}, OUT_12_14);
	wire [3:0] OUT_12_15;
	CAS CAS_12_15( {OUT_12_14[0], OUT_11_14[1], M[15], Q[20]}, OUT_12_15);
	wire [3:0] OUT_12_16;
	CAS CAS_12_16( {OUT_12_15[0], OUT_11_15[1], M[16], Q[20]}, OUT_12_16);
	wire [3:0] OUT_12_17;
	CAS CAS_12_17( {OUT_12_16[0], OUT_11_16[1], M[17], Q[20]}, OUT_12_17);
	wire [3:0] OUT_12_18;
	CAS CAS_12_18( {OUT_12_17[0], OUT_11_17[1], M[18], Q[20]}, OUT_12_18);
	wire [3:0] OUT_12_19;
	CAS CAS_12_19( {OUT_12_18[0], OUT_11_18[1], M[19], Q[20]}, OUT_12_19);
	wire [3:0] OUT_12_20;
	CAS CAS_12_20( {OUT_12_19[0], OUT_11_19[1], M[20], Q[20]}, OUT_12_20);
	wire [3:0] OUT_12_21;
	CAS CAS_12_21( {OUT_12_20[0], OUT_11_20[1], M[21], Q[20]}, OUT_12_21);
	wire [3:0] OUT_12_22;
	CAS CAS_12_22( {OUT_12_21[0], OUT_11_21[1], M[22], Q[20]}, OUT_12_22);
	wire [3:0] OUT_12_23;
	CAS CAS_12_23( {OUT_12_22[0], OUT_11_22[1], M[23], Q[20]}, OUT_12_23);
	wire [3:0] OUT_12_24;
	CAS CAS_12_24( {OUT_12_23[0], OUT_11_23[1], M[24], Q[20]}, OUT_12_24);
	wire [3:0] OUT_12_25;
	CAS CAS_12_25( {OUT_12_24[0], OUT_11_24[1], M[25], Q[20]}, OUT_12_25);
	wire [3:0] OUT_12_26;
	CAS CAS_12_26( {OUT_12_25[0], OUT_11_25[1], M[26], Q[20]}, OUT_12_26);
	wire [3:0] OUT_12_27;
	CAS CAS_12_27( {OUT_12_26[0], OUT_11_26[1], M[27], Q[20]}, OUT_12_27);
	wire [3:0] OUT_12_28;
	CAS CAS_12_28( {OUT_12_27[0], OUT_11_27[1], M[28], Q[20]}, OUT_12_28);
	wire [3:0] OUT_12_29;
	CAS CAS_12_29( {OUT_12_28[0], OUT_11_28[1], M[29], Q[20]}, OUT_12_29);
	wire [3:0] OUT_12_30;
	CAS CAS_12_30( {OUT_12_29[0], OUT_11_29[1], M[30], Q[20]}, OUT_12_30);
	wire [3:0] OUT_12_31;
	CAS CAS_12_31( {OUT_12_30[0], OUT_11_30[1], M[31], Q[20]}, OUT_12_31);
	assign Q[19] = OUT_12_31[0];

// Level - 14
	wire [3:0] OUT_13_0;
	CAS CAS_13_0( {Q[19], D[18], M[0], Q[19]}, OUT_13_0);
	wire [3:0] OUT_13_1;
	CAS CAS_13_1( {OUT_13_0[0], OUT_12_0[1], M[1], Q[19]}, OUT_13_1);
	wire [3:0] OUT_13_2;
	CAS CAS_13_2( {OUT_13_1[0], OUT_12_1[1], M[2], Q[19]}, OUT_13_2);
	wire [3:0] OUT_13_3;
	CAS CAS_13_3( {OUT_13_2[0], OUT_12_2[1], M[3], Q[19]}, OUT_13_3);
	wire [3:0] OUT_13_4;
	CAS CAS_13_4( {OUT_13_3[0], OUT_12_3[1], M[4], Q[19]}, OUT_13_4);
	wire [3:0] OUT_13_5;
	CAS CAS_13_5( {OUT_13_4[0], OUT_12_4[1], M[5], Q[19]}, OUT_13_5);
	wire [3:0] OUT_13_6;
	CAS CAS_13_6( {OUT_13_5[0], OUT_12_5[1], M[6], Q[19]}, OUT_13_6);
	wire [3:0] OUT_13_7;
	CAS CAS_13_7( {OUT_13_6[0], OUT_12_6[1], M[7], Q[19]}, OUT_13_7);
	wire [3:0] OUT_13_8;
	CAS CAS_13_8( {OUT_13_7[0], OUT_12_7[1], M[8], Q[19]}, OUT_13_8);
	wire [3:0] OUT_13_9;
	CAS CAS_13_9( {OUT_13_8[0], OUT_12_8[1], M[9], Q[19]}, OUT_13_9);
	wire [3:0] OUT_13_10;
	CAS CAS_13_10( {OUT_13_9[0], OUT_12_9[1], M[10], Q[19]}, OUT_13_10);
	wire [3:0] OUT_13_11;
	CAS CAS_13_11( {OUT_13_10[0], OUT_12_10[1], M[11], Q[19]}, OUT_13_11);
	wire [3:0] OUT_13_12;
	CAS CAS_13_12( {OUT_13_11[0], OUT_12_11[1], M[12], Q[19]}, OUT_13_12);
	wire [3:0] OUT_13_13;
	CAS CAS_13_13( {OUT_13_12[0], OUT_12_12[1], M[13], Q[19]}, OUT_13_13);
	wire [3:0] OUT_13_14;
	CAS CAS_13_14( {OUT_13_13[0], OUT_12_13[1], M[14], Q[19]}, OUT_13_14);
	wire [3:0] OUT_13_15;
	CAS CAS_13_15( {OUT_13_14[0], OUT_12_14[1], M[15], Q[19]}, OUT_13_15);
	wire [3:0] OUT_13_16;
	CAS CAS_13_16( {OUT_13_15[0], OUT_12_15[1], M[16], Q[19]}, OUT_13_16);
	wire [3:0] OUT_13_17;
	CAS CAS_13_17( {OUT_13_16[0], OUT_12_16[1], M[17], Q[19]}, OUT_13_17);
	wire [3:0] OUT_13_18;
	CAS CAS_13_18( {OUT_13_17[0], OUT_12_17[1], M[18], Q[19]}, OUT_13_18);
	wire [3:0] OUT_13_19;
	CAS CAS_13_19( {OUT_13_18[0], OUT_12_18[1], M[19], Q[19]}, OUT_13_19);
	wire [3:0] OUT_13_20;
	CAS CAS_13_20( {OUT_13_19[0], OUT_12_19[1], M[20], Q[19]}, OUT_13_20);
	wire [3:0] OUT_13_21;
	CAS CAS_13_21( {OUT_13_20[0], OUT_12_20[1], M[21], Q[19]}, OUT_13_21);
	wire [3:0] OUT_13_22;
	CAS CAS_13_22( {OUT_13_21[0], OUT_12_21[1], M[22], Q[19]}, OUT_13_22);
	wire [3:0] OUT_13_23;
	CAS CAS_13_23( {OUT_13_22[0], OUT_12_22[1], M[23], Q[19]}, OUT_13_23);
	wire [3:0] OUT_13_24;
	CAS CAS_13_24( {OUT_13_23[0], OUT_12_23[1], M[24], Q[19]}, OUT_13_24);
	wire [3:0] OUT_13_25;
	CAS CAS_13_25( {OUT_13_24[0], OUT_12_24[1], M[25], Q[19]}, OUT_13_25);
	wire [3:0] OUT_13_26;
	CAS CAS_13_26( {OUT_13_25[0], OUT_12_25[1], M[26], Q[19]}, OUT_13_26);
	wire [3:0] OUT_13_27;
	CAS CAS_13_27( {OUT_13_26[0], OUT_12_26[1], M[27], Q[19]}, OUT_13_27);
	wire [3:0] OUT_13_28;
	CAS CAS_13_28( {OUT_13_27[0], OUT_12_27[1], M[28], Q[19]}, OUT_13_28);
	wire [3:0] OUT_13_29;
	CAS CAS_13_29( {OUT_13_28[0], OUT_12_28[1], M[29], Q[19]}, OUT_13_29);
	wire [3:0] OUT_13_30;
	CAS CAS_13_30( {OUT_13_29[0], OUT_12_29[1], M[30], Q[19]}, OUT_13_30);
	wire [3:0] OUT_13_31;
	CAS CAS_13_31( {OUT_13_30[0], OUT_12_30[1], M[31], Q[19]}, OUT_13_31);
	assign Q[18] = OUT_13_31[0];

// Level - 15
	wire [3:0] OUT_14_0;
	CAS CAS_14_0( {Q[18], D[17], M[0], Q[18]}, OUT_14_0);
	wire [3:0] OUT_14_1;
	CAS CAS_14_1( {OUT_14_0[0], OUT_13_0[1], M[1], Q[18]}, OUT_14_1);
	wire [3:0] OUT_14_2;
	CAS CAS_14_2( {OUT_14_1[0], OUT_13_1[1], M[2], Q[18]}, OUT_14_2);
	wire [3:0] OUT_14_3;
	CAS CAS_14_3( {OUT_14_2[0], OUT_13_2[1], M[3], Q[18]}, OUT_14_3);
	wire [3:0] OUT_14_4;
	CAS CAS_14_4( {OUT_14_3[0], OUT_13_3[1], M[4], Q[18]}, OUT_14_4);
	wire [3:0] OUT_14_5;
	CAS CAS_14_5( {OUT_14_4[0], OUT_13_4[1], M[5], Q[18]}, OUT_14_5);
	wire [3:0] OUT_14_6;
	CAS CAS_14_6( {OUT_14_5[0], OUT_13_5[1], M[6], Q[18]}, OUT_14_6);
	wire [3:0] OUT_14_7;
	CAS CAS_14_7( {OUT_14_6[0], OUT_13_6[1], M[7], Q[18]}, OUT_14_7);
	wire [3:0] OUT_14_8;
	CAS CAS_14_8( {OUT_14_7[0], OUT_13_7[1], M[8], Q[18]}, OUT_14_8);
	wire [3:0] OUT_14_9;
	CAS CAS_14_9( {OUT_14_8[0], OUT_13_8[1], M[9], Q[18]}, OUT_14_9);
	wire [3:0] OUT_14_10;
	CAS CAS_14_10( {OUT_14_9[0], OUT_13_9[1], M[10], Q[18]}, OUT_14_10);
	wire [3:0] OUT_14_11;
	CAS CAS_14_11( {OUT_14_10[0], OUT_13_10[1], M[11], Q[18]}, OUT_14_11);
	wire [3:0] OUT_14_12;
	CAS CAS_14_12( {OUT_14_11[0], OUT_13_11[1], M[12], Q[18]}, OUT_14_12);
	wire [3:0] OUT_14_13;
	CAS CAS_14_13( {OUT_14_12[0], OUT_13_12[1], M[13], Q[18]}, OUT_14_13);
	wire [3:0] OUT_14_14;
	CAS CAS_14_14( {OUT_14_13[0], OUT_13_13[1], M[14], Q[18]}, OUT_14_14);
	wire [3:0] OUT_14_15;
	CAS CAS_14_15( {OUT_14_14[0], OUT_13_14[1], M[15], Q[18]}, OUT_14_15);
	wire [3:0] OUT_14_16;
	CAS CAS_14_16( {OUT_14_15[0], OUT_13_15[1], M[16], Q[18]}, OUT_14_16);
	wire [3:0] OUT_14_17;
	CAS CAS_14_17( {OUT_14_16[0], OUT_13_16[1], M[17], Q[18]}, OUT_14_17);
	wire [3:0] OUT_14_18;
	CAS CAS_14_18( {OUT_14_17[0], OUT_13_17[1], M[18], Q[18]}, OUT_14_18);
	wire [3:0] OUT_14_19;
	CAS CAS_14_19( {OUT_14_18[0], OUT_13_18[1], M[19], Q[18]}, OUT_14_19);
	wire [3:0] OUT_14_20;
	CAS CAS_14_20( {OUT_14_19[0], OUT_13_19[1], M[20], Q[18]}, OUT_14_20);
	wire [3:0] OUT_14_21;
	CAS CAS_14_21( {OUT_14_20[0], OUT_13_20[1], M[21], Q[18]}, OUT_14_21);
	wire [3:0] OUT_14_22;
	CAS CAS_14_22( {OUT_14_21[0], OUT_13_21[1], M[22], Q[18]}, OUT_14_22);
	wire [3:0] OUT_14_23;
	CAS CAS_14_23( {OUT_14_22[0], OUT_13_22[1], M[23], Q[18]}, OUT_14_23);
	wire [3:0] OUT_14_24;
	CAS CAS_14_24( {OUT_14_23[0], OUT_13_23[1], M[24], Q[18]}, OUT_14_24);
	wire [3:0] OUT_14_25;
	CAS CAS_14_25( {OUT_14_24[0], OUT_13_24[1], M[25], Q[18]}, OUT_14_25);
	wire [3:0] OUT_14_26;
	CAS CAS_14_26( {OUT_14_25[0], OUT_13_25[1], M[26], Q[18]}, OUT_14_26);
	wire [3:0] OUT_14_27;
	CAS CAS_14_27( {OUT_14_26[0], OUT_13_26[1], M[27], Q[18]}, OUT_14_27);
	wire [3:0] OUT_14_28;
	CAS CAS_14_28( {OUT_14_27[0], OUT_13_27[1], M[28], Q[18]}, OUT_14_28);
	wire [3:0] OUT_14_29;
	CAS CAS_14_29( {OUT_14_28[0], OUT_13_28[1], M[29], Q[18]}, OUT_14_29);
	wire [3:0] OUT_14_30;
	CAS CAS_14_30( {OUT_14_29[0], OUT_13_29[1], M[30], Q[18]}, OUT_14_30);
	wire [3:0] OUT_14_31;
	CAS CAS_14_31( {OUT_14_30[0], OUT_13_30[1], M[31], Q[18]}, OUT_14_31);
	assign Q[17] = OUT_14_31[0];

// Level - 16
	wire [3:0] OUT_15_0;
	CAS CAS_15_0( {Q[17], D[16], M[0], Q[17]}, OUT_15_0);
	wire [3:0] OUT_15_1;
	CAS CAS_15_1( {OUT_15_0[0], OUT_14_0[1], M[1], Q[17]}, OUT_15_1);
	wire [3:0] OUT_15_2;
	CAS CAS_15_2( {OUT_15_1[0], OUT_14_1[1], M[2], Q[17]}, OUT_15_2);
	wire [3:0] OUT_15_3;
	CAS CAS_15_3( {OUT_15_2[0], OUT_14_2[1], M[3], Q[17]}, OUT_15_3);
	wire [3:0] OUT_15_4;
	CAS CAS_15_4( {OUT_15_3[0], OUT_14_3[1], M[4], Q[17]}, OUT_15_4);
	wire [3:0] OUT_15_5;
	CAS CAS_15_5( {OUT_15_4[0], OUT_14_4[1], M[5], Q[17]}, OUT_15_5);
	wire [3:0] OUT_15_6;
	CAS CAS_15_6( {OUT_15_5[0], OUT_14_5[1], M[6], Q[17]}, OUT_15_6);
	wire [3:0] OUT_15_7;
	CAS CAS_15_7( {OUT_15_6[0], OUT_14_6[1], M[7], Q[17]}, OUT_15_7);
	wire [3:0] OUT_15_8;
	CAS CAS_15_8( {OUT_15_7[0], OUT_14_7[1], M[8], Q[17]}, OUT_15_8);
	wire [3:0] OUT_15_9;
	CAS CAS_15_9( {OUT_15_8[0], OUT_14_8[1], M[9], Q[17]}, OUT_15_9);
	wire [3:0] OUT_15_10;
	CAS CAS_15_10( {OUT_15_9[0], OUT_14_9[1], M[10], Q[17]}, OUT_15_10);
	wire [3:0] OUT_15_11;
	CAS CAS_15_11( {OUT_15_10[0], OUT_14_10[1], M[11], Q[17]}, OUT_15_11);
	wire [3:0] OUT_15_12;
	CAS CAS_15_12( {OUT_15_11[0], OUT_14_11[1], M[12], Q[17]}, OUT_15_12);
	wire [3:0] OUT_15_13;
	CAS CAS_15_13( {OUT_15_12[0], OUT_14_12[1], M[13], Q[17]}, OUT_15_13);
	wire [3:0] OUT_15_14;
	CAS CAS_15_14( {OUT_15_13[0], OUT_14_13[1], M[14], Q[17]}, OUT_15_14);
	wire [3:0] OUT_15_15;
	CAS CAS_15_15( {OUT_15_14[0], OUT_14_14[1], M[15], Q[17]}, OUT_15_15);
	wire [3:0] OUT_15_16;
	CAS CAS_15_16( {OUT_15_15[0], OUT_14_15[1], M[16], Q[17]}, OUT_15_16);
	wire [3:0] OUT_15_17;
	CAS CAS_15_17( {OUT_15_16[0], OUT_14_16[1], M[17], Q[17]}, OUT_15_17);
	wire [3:0] OUT_15_18;
	CAS CAS_15_18( {OUT_15_17[0], OUT_14_17[1], M[18], Q[17]}, OUT_15_18);
	wire [3:0] OUT_15_19;
	CAS CAS_15_19( {OUT_15_18[0], OUT_14_18[1], M[19], Q[17]}, OUT_15_19);
	wire [3:0] OUT_15_20;
	CAS CAS_15_20( {OUT_15_19[0], OUT_14_19[1], M[20], Q[17]}, OUT_15_20);
	wire [3:0] OUT_15_21;
	CAS CAS_15_21( {OUT_15_20[0], OUT_14_20[1], M[21], Q[17]}, OUT_15_21);
	wire [3:0] OUT_15_22;
	CAS CAS_15_22( {OUT_15_21[0], OUT_14_21[1], M[22], Q[17]}, OUT_15_22);
	wire [3:0] OUT_15_23;
	CAS CAS_15_23( {OUT_15_22[0], OUT_14_22[1], M[23], Q[17]}, OUT_15_23);
	wire [3:0] OUT_15_24;
	CAS CAS_15_24( {OUT_15_23[0], OUT_14_23[1], M[24], Q[17]}, OUT_15_24);
	wire [3:0] OUT_15_25;
	CAS CAS_15_25( {OUT_15_24[0], OUT_14_24[1], M[25], Q[17]}, OUT_15_25);
	wire [3:0] OUT_15_26;
	CAS CAS_15_26( {OUT_15_25[0], OUT_14_25[1], M[26], Q[17]}, OUT_15_26);
	wire [3:0] OUT_15_27;
	CAS CAS_15_27( {OUT_15_26[0], OUT_14_26[1], M[27], Q[17]}, OUT_15_27);
	wire [3:0] OUT_15_28;
	CAS CAS_15_28( {OUT_15_27[0], OUT_14_27[1], M[28], Q[17]}, OUT_15_28);
	wire [3:0] OUT_15_29;
	CAS CAS_15_29( {OUT_15_28[0], OUT_14_28[1], M[29], Q[17]}, OUT_15_29);
	wire [3:0] OUT_15_30;
	CAS CAS_15_30( {OUT_15_29[0], OUT_14_29[1], M[30], Q[17]}, OUT_15_30);
	wire [3:0] OUT_15_31;
	CAS CAS_15_31( {OUT_15_30[0], OUT_14_30[1], M[31], Q[17]}, OUT_15_31);
	assign Q[16] = OUT_15_31[0];

// Level - 17
	wire [3:0] OUT_16_0;
	CAS CAS_16_0( {Q[16], D[15], M[0], Q[16]}, OUT_16_0);
	wire [3:0] OUT_16_1;
	CAS CAS_16_1( {OUT_16_0[0], OUT_15_0[1], M[1], Q[16]}, OUT_16_1);
	wire [3:0] OUT_16_2;
	CAS CAS_16_2( {OUT_16_1[0], OUT_15_1[1], M[2], Q[16]}, OUT_16_2);
	wire [3:0] OUT_16_3;
	CAS CAS_16_3( {OUT_16_2[0], OUT_15_2[1], M[3], Q[16]}, OUT_16_3);
	wire [3:0] OUT_16_4;
	CAS CAS_16_4( {OUT_16_3[0], OUT_15_3[1], M[4], Q[16]}, OUT_16_4);
	wire [3:0] OUT_16_5;
	CAS CAS_16_5( {OUT_16_4[0], OUT_15_4[1], M[5], Q[16]}, OUT_16_5);
	wire [3:0] OUT_16_6;
	CAS CAS_16_6( {OUT_16_5[0], OUT_15_5[1], M[6], Q[16]}, OUT_16_6);
	wire [3:0] OUT_16_7;
	CAS CAS_16_7( {OUT_16_6[0], OUT_15_6[1], M[7], Q[16]}, OUT_16_7);
	wire [3:0] OUT_16_8;
	CAS CAS_16_8( {OUT_16_7[0], OUT_15_7[1], M[8], Q[16]}, OUT_16_8);
	wire [3:0] OUT_16_9;
	CAS CAS_16_9( {OUT_16_8[0], OUT_15_8[1], M[9], Q[16]}, OUT_16_9);
	wire [3:0] OUT_16_10;
	CAS CAS_16_10( {OUT_16_9[0], OUT_15_9[1], M[10], Q[16]}, OUT_16_10);
	wire [3:0] OUT_16_11;
	CAS CAS_16_11( {OUT_16_10[0], OUT_15_10[1], M[11], Q[16]}, OUT_16_11);
	wire [3:0] OUT_16_12;
	CAS CAS_16_12( {OUT_16_11[0], OUT_15_11[1], M[12], Q[16]}, OUT_16_12);
	wire [3:0] OUT_16_13;
	CAS CAS_16_13( {OUT_16_12[0], OUT_15_12[1], M[13], Q[16]}, OUT_16_13);
	wire [3:0] OUT_16_14;
	CAS CAS_16_14( {OUT_16_13[0], OUT_15_13[1], M[14], Q[16]}, OUT_16_14);
	wire [3:0] OUT_16_15;
	CAS CAS_16_15( {OUT_16_14[0], OUT_15_14[1], M[15], Q[16]}, OUT_16_15);
	wire [3:0] OUT_16_16;
	CAS CAS_16_16( {OUT_16_15[0], OUT_15_15[1], M[16], Q[16]}, OUT_16_16);
	wire [3:0] OUT_16_17;
	CAS CAS_16_17( {OUT_16_16[0], OUT_15_16[1], M[17], Q[16]}, OUT_16_17);
	wire [3:0] OUT_16_18;
	CAS CAS_16_18( {OUT_16_17[0], OUT_15_17[1], M[18], Q[16]}, OUT_16_18);
	wire [3:0] OUT_16_19;
	CAS CAS_16_19( {OUT_16_18[0], OUT_15_18[1], M[19], Q[16]}, OUT_16_19);
	wire [3:0] OUT_16_20;
	CAS CAS_16_20( {OUT_16_19[0], OUT_15_19[1], M[20], Q[16]}, OUT_16_20);
	wire [3:0] OUT_16_21;
	CAS CAS_16_21( {OUT_16_20[0], OUT_15_20[1], M[21], Q[16]}, OUT_16_21);
	wire [3:0] OUT_16_22;
	CAS CAS_16_22( {OUT_16_21[0], OUT_15_21[1], M[22], Q[16]}, OUT_16_22);
	wire [3:0] OUT_16_23;
	CAS CAS_16_23( {OUT_16_22[0], OUT_15_22[1], M[23], Q[16]}, OUT_16_23);
	wire [3:0] OUT_16_24;
	CAS CAS_16_24( {OUT_16_23[0], OUT_15_23[1], M[24], Q[16]}, OUT_16_24);
	wire [3:0] OUT_16_25;
	CAS CAS_16_25( {OUT_16_24[0], OUT_15_24[1], M[25], Q[16]}, OUT_16_25);
	wire [3:0] OUT_16_26;
	CAS CAS_16_26( {OUT_16_25[0], OUT_15_25[1], M[26], Q[16]}, OUT_16_26);
	wire [3:0] OUT_16_27;
	CAS CAS_16_27( {OUT_16_26[0], OUT_15_26[1], M[27], Q[16]}, OUT_16_27);
	wire [3:0] OUT_16_28;
	CAS CAS_16_28( {OUT_16_27[0], OUT_15_27[1], M[28], Q[16]}, OUT_16_28);
	wire [3:0] OUT_16_29;
	CAS CAS_16_29( {OUT_16_28[0], OUT_15_28[1], M[29], Q[16]}, OUT_16_29);
	wire [3:0] OUT_16_30;
	CAS CAS_16_30( {OUT_16_29[0], OUT_15_29[1], M[30], Q[16]}, OUT_16_30);
	wire [3:0] OUT_16_31;
	CAS CAS_16_31( {OUT_16_30[0], OUT_15_30[1], M[31], Q[16]}, OUT_16_31);
	assign Q[15] = OUT_16_31[0];

// Level - 18
	wire [3:0] OUT_17_0;
	CAS CAS_17_0( {Q[15], D[14], M[0], Q[15]}, OUT_17_0);
	wire [3:0] OUT_17_1;
	CAS CAS_17_1( {OUT_17_0[0], OUT_16_0[1], M[1], Q[15]}, OUT_17_1);
	wire [3:0] OUT_17_2;
	CAS CAS_17_2( {OUT_17_1[0], OUT_16_1[1], M[2], Q[15]}, OUT_17_2);
	wire [3:0] OUT_17_3;
	CAS CAS_17_3( {OUT_17_2[0], OUT_16_2[1], M[3], Q[15]}, OUT_17_3);
	wire [3:0] OUT_17_4;
	CAS CAS_17_4( {OUT_17_3[0], OUT_16_3[1], M[4], Q[15]}, OUT_17_4);
	wire [3:0] OUT_17_5;
	CAS CAS_17_5( {OUT_17_4[0], OUT_16_4[1], M[5], Q[15]}, OUT_17_5);
	wire [3:0] OUT_17_6;
	CAS CAS_17_6( {OUT_17_5[0], OUT_16_5[1], M[6], Q[15]}, OUT_17_6);
	wire [3:0] OUT_17_7;
	CAS CAS_17_7( {OUT_17_6[0], OUT_16_6[1], M[7], Q[15]}, OUT_17_7);
	wire [3:0] OUT_17_8;
	CAS CAS_17_8( {OUT_17_7[0], OUT_16_7[1], M[8], Q[15]}, OUT_17_8);
	wire [3:0] OUT_17_9;
	CAS CAS_17_9( {OUT_17_8[0], OUT_16_8[1], M[9], Q[15]}, OUT_17_9);
	wire [3:0] OUT_17_10;
	CAS CAS_17_10( {OUT_17_9[0], OUT_16_9[1], M[10], Q[15]}, OUT_17_10);
	wire [3:0] OUT_17_11;
	CAS CAS_17_11( {OUT_17_10[0], OUT_16_10[1], M[11], Q[15]}, OUT_17_11);
	wire [3:0] OUT_17_12;
	CAS CAS_17_12( {OUT_17_11[0], OUT_16_11[1], M[12], Q[15]}, OUT_17_12);
	wire [3:0] OUT_17_13;
	CAS CAS_17_13( {OUT_17_12[0], OUT_16_12[1], M[13], Q[15]}, OUT_17_13);
	wire [3:0] OUT_17_14;
	CAS CAS_17_14( {OUT_17_13[0], OUT_16_13[1], M[14], Q[15]}, OUT_17_14);
	wire [3:0] OUT_17_15;
	CAS CAS_17_15( {OUT_17_14[0], OUT_16_14[1], M[15], Q[15]}, OUT_17_15);
	wire [3:0] OUT_17_16;
	CAS CAS_17_16( {OUT_17_15[0], OUT_16_15[1], M[16], Q[15]}, OUT_17_16);
	wire [3:0] OUT_17_17;
	CAS CAS_17_17( {OUT_17_16[0], OUT_16_16[1], M[17], Q[15]}, OUT_17_17);
	wire [3:0] OUT_17_18;
	CAS CAS_17_18( {OUT_17_17[0], OUT_16_17[1], M[18], Q[15]}, OUT_17_18);
	wire [3:0] OUT_17_19;
	CAS CAS_17_19( {OUT_17_18[0], OUT_16_18[1], M[19], Q[15]}, OUT_17_19);
	wire [3:0] OUT_17_20;
	CAS CAS_17_20( {OUT_17_19[0], OUT_16_19[1], M[20], Q[15]}, OUT_17_20);
	wire [3:0] OUT_17_21;
	CAS CAS_17_21( {OUT_17_20[0], OUT_16_20[1], M[21], Q[15]}, OUT_17_21);
	wire [3:0] OUT_17_22;
	CAS CAS_17_22( {OUT_17_21[0], OUT_16_21[1], M[22], Q[15]}, OUT_17_22);
	wire [3:0] OUT_17_23;
	CAS CAS_17_23( {OUT_17_22[0], OUT_16_22[1], M[23], Q[15]}, OUT_17_23);
	wire [3:0] OUT_17_24;
	CAS CAS_17_24( {OUT_17_23[0], OUT_16_23[1], M[24], Q[15]}, OUT_17_24);
	wire [3:0] OUT_17_25;
	CAS CAS_17_25( {OUT_17_24[0], OUT_16_24[1], M[25], Q[15]}, OUT_17_25);
	wire [3:0] OUT_17_26;
	CAS CAS_17_26( {OUT_17_25[0], OUT_16_25[1], M[26], Q[15]}, OUT_17_26);
	wire [3:0] OUT_17_27;
	CAS CAS_17_27( {OUT_17_26[0], OUT_16_26[1], M[27], Q[15]}, OUT_17_27);
	wire [3:0] OUT_17_28;
	CAS CAS_17_28( {OUT_17_27[0], OUT_16_27[1], M[28], Q[15]}, OUT_17_28);
	wire [3:0] OUT_17_29;
	CAS CAS_17_29( {OUT_17_28[0], OUT_16_28[1], M[29], Q[15]}, OUT_17_29);
	wire [3:0] OUT_17_30;
	CAS CAS_17_30( {OUT_17_29[0], OUT_16_29[1], M[30], Q[15]}, OUT_17_30);
	wire [3:0] OUT_17_31;
	CAS CAS_17_31( {OUT_17_30[0], OUT_16_30[1], M[31], Q[15]}, OUT_17_31);
	assign Q[14] = OUT_17_31[0];

// Level - 19
	wire [3:0] OUT_18_0;
	CAS CAS_18_0( {Q[14], D[13], M[0], Q[14]}, OUT_18_0);
	wire [3:0] OUT_18_1;
	CAS CAS_18_1( {OUT_18_0[0], OUT_17_0[1], M[1], Q[14]}, OUT_18_1);
	wire [3:0] OUT_18_2;
	CAS CAS_18_2( {OUT_18_1[0], OUT_17_1[1], M[2], Q[14]}, OUT_18_2);
	wire [3:0] OUT_18_3;
	CAS CAS_18_3( {OUT_18_2[0], OUT_17_2[1], M[3], Q[14]}, OUT_18_3);
	wire [3:0] OUT_18_4;
	CAS CAS_18_4( {OUT_18_3[0], OUT_17_3[1], M[4], Q[14]}, OUT_18_4);
	wire [3:0] OUT_18_5;
	CAS CAS_18_5( {OUT_18_4[0], OUT_17_4[1], M[5], Q[14]}, OUT_18_5);
	wire [3:0] OUT_18_6;
	CAS CAS_18_6( {OUT_18_5[0], OUT_17_5[1], M[6], Q[14]}, OUT_18_6);
	wire [3:0] OUT_18_7;
	CAS CAS_18_7( {OUT_18_6[0], OUT_17_6[1], M[7], Q[14]}, OUT_18_7);
	wire [3:0] OUT_18_8;
	CAS CAS_18_8( {OUT_18_7[0], OUT_17_7[1], M[8], Q[14]}, OUT_18_8);
	wire [3:0] OUT_18_9;
	CAS CAS_18_9( {OUT_18_8[0], OUT_17_8[1], M[9], Q[14]}, OUT_18_9);
	wire [3:0] OUT_18_10;
	CAS CAS_18_10( {OUT_18_9[0], OUT_17_9[1], M[10], Q[14]}, OUT_18_10);
	wire [3:0] OUT_18_11;
	CAS CAS_18_11( {OUT_18_10[0], OUT_17_10[1], M[11], Q[14]}, OUT_18_11);
	wire [3:0] OUT_18_12;
	CAS CAS_18_12( {OUT_18_11[0], OUT_17_11[1], M[12], Q[14]}, OUT_18_12);
	wire [3:0] OUT_18_13;
	CAS CAS_18_13( {OUT_18_12[0], OUT_17_12[1], M[13], Q[14]}, OUT_18_13);
	wire [3:0] OUT_18_14;
	CAS CAS_18_14( {OUT_18_13[0], OUT_17_13[1], M[14], Q[14]}, OUT_18_14);
	wire [3:0] OUT_18_15;
	CAS CAS_18_15( {OUT_18_14[0], OUT_17_14[1], M[15], Q[14]}, OUT_18_15);
	wire [3:0] OUT_18_16;
	CAS CAS_18_16( {OUT_18_15[0], OUT_17_15[1], M[16], Q[14]}, OUT_18_16);
	wire [3:0] OUT_18_17;
	CAS CAS_18_17( {OUT_18_16[0], OUT_17_16[1], M[17], Q[14]}, OUT_18_17);
	wire [3:0] OUT_18_18;
	CAS CAS_18_18( {OUT_18_17[0], OUT_17_17[1], M[18], Q[14]}, OUT_18_18);
	wire [3:0] OUT_18_19;
	CAS CAS_18_19( {OUT_18_18[0], OUT_17_18[1], M[19], Q[14]}, OUT_18_19);
	wire [3:0] OUT_18_20;
	CAS CAS_18_20( {OUT_18_19[0], OUT_17_19[1], M[20], Q[14]}, OUT_18_20);
	wire [3:0] OUT_18_21;
	CAS CAS_18_21( {OUT_18_20[0], OUT_17_20[1], M[21], Q[14]}, OUT_18_21);
	wire [3:0] OUT_18_22;
	CAS CAS_18_22( {OUT_18_21[0], OUT_17_21[1], M[22], Q[14]}, OUT_18_22);
	wire [3:0] OUT_18_23;
	CAS CAS_18_23( {OUT_18_22[0], OUT_17_22[1], M[23], Q[14]}, OUT_18_23);
	wire [3:0] OUT_18_24;
	CAS CAS_18_24( {OUT_18_23[0], OUT_17_23[1], M[24], Q[14]}, OUT_18_24);
	wire [3:0] OUT_18_25;
	CAS CAS_18_25( {OUT_18_24[0], OUT_17_24[1], M[25], Q[14]}, OUT_18_25);
	wire [3:0] OUT_18_26;
	CAS CAS_18_26( {OUT_18_25[0], OUT_17_25[1], M[26], Q[14]}, OUT_18_26);
	wire [3:0] OUT_18_27;
	CAS CAS_18_27( {OUT_18_26[0], OUT_17_26[1], M[27], Q[14]}, OUT_18_27);
	wire [3:0] OUT_18_28;
	CAS CAS_18_28( {OUT_18_27[0], OUT_17_27[1], M[28], Q[14]}, OUT_18_28);
	wire [3:0] OUT_18_29;
	CAS CAS_18_29( {OUT_18_28[0], OUT_17_28[1], M[29], Q[14]}, OUT_18_29);
	wire [3:0] OUT_18_30;
	CAS CAS_18_30( {OUT_18_29[0], OUT_17_29[1], M[30], Q[14]}, OUT_18_30);
	wire [3:0] OUT_18_31;
	CAS CAS_18_31( {OUT_18_30[0], OUT_17_30[1], M[31], Q[14]}, OUT_18_31);
	assign Q[13] = OUT_18_31[0];

// Level - 20
	wire [3:0] OUT_19_0;
	CAS CAS_19_0( {Q[13], D[12], M[0], Q[13]}, OUT_19_0);
	wire [3:0] OUT_19_1;
	CAS CAS_19_1( {OUT_19_0[0], OUT_18_0[1], M[1], Q[13]}, OUT_19_1);
	wire [3:0] OUT_19_2;
	CAS CAS_19_2( {OUT_19_1[0], OUT_18_1[1], M[2], Q[13]}, OUT_19_2);
	wire [3:0] OUT_19_3;
	CAS CAS_19_3( {OUT_19_2[0], OUT_18_2[1], M[3], Q[13]}, OUT_19_3);
	wire [3:0] OUT_19_4;
	CAS CAS_19_4( {OUT_19_3[0], OUT_18_3[1], M[4], Q[13]}, OUT_19_4);
	wire [3:0] OUT_19_5;
	CAS CAS_19_5( {OUT_19_4[0], OUT_18_4[1], M[5], Q[13]}, OUT_19_5);
	wire [3:0] OUT_19_6;
	CAS CAS_19_6( {OUT_19_5[0], OUT_18_5[1], M[6], Q[13]}, OUT_19_6);
	wire [3:0] OUT_19_7;
	CAS CAS_19_7( {OUT_19_6[0], OUT_18_6[1], M[7], Q[13]}, OUT_19_7);
	wire [3:0] OUT_19_8;
	CAS CAS_19_8( {OUT_19_7[0], OUT_18_7[1], M[8], Q[13]}, OUT_19_8);
	wire [3:0] OUT_19_9;
	CAS CAS_19_9( {OUT_19_8[0], OUT_18_8[1], M[9], Q[13]}, OUT_19_9);
	wire [3:0] OUT_19_10;
	CAS CAS_19_10( {OUT_19_9[0], OUT_18_9[1], M[10], Q[13]}, OUT_19_10);
	wire [3:0] OUT_19_11;
	CAS CAS_19_11( {OUT_19_10[0], OUT_18_10[1], M[11], Q[13]}, OUT_19_11);
	wire [3:0] OUT_19_12;
	CAS CAS_19_12( {OUT_19_11[0], OUT_18_11[1], M[12], Q[13]}, OUT_19_12);
	wire [3:0] OUT_19_13;
	CAS CAS_19_13( {OUT_19_12[0], OUT_18_12[1], M[13], Q[13]}, OUT_19_13);
	wire [3:0] OUT_19_14;
	CAS CAS_19_14( {OUT_19_13[0], OUT_18_13[1], M[14], Q[13]}, OUT_19_14);
	wire [3:0] OUT_19_15;
	CAS CAS_19_15( {OUT_19_14[0], OUT_18_14[1], M[15], Q[13]}, OUT_19_15);
	wire [3:0] OUT_19_16;
	CAS CAS_19_16( {OUT_19_15[0], OUT_18_15[1], M[16], Q[13]}, OUT_19_16);
	wire [3:0] OUT_19_17;
	CAS CAS_19_17( {OUT_19_16[0], OUT_18_16[1], M[17], Q[13]}, OUT_19_17);
	wire [3:0] OUT_19_18;
	CAS CAS_19_18( {OUT_19_17[0], OUT_18_17[1], M[18], Q[13]}, OUT_19_18);
	wire [3:0] OUT_19_19;
	CAS CAS_19_19( {OUT_19_18[0], OUT_18_18[1], M[19], Q[13]}, OUT_19_19);
	wire [3:0] OUT_19_20;
	CAS CAS_19_20( {OUT_19_19[0], OUT_18_19[1], M[20], Q[13]}, OUT_19_20);
	wire [3:0] OUT_19_21;
	CAS CAS_19_21( {OUT_19_20[0], OUT_18_20[1], M[21], Q[13]}, OUT_19_21);
	wire [3:0] OUT_19_22;
	CAS CAS_19_22( {OUT_19_21[0], OUT_18_21[1], M[22], Q[13]}, OUT_19_22);
	wire [3:0] OUT_19_23;
	CAS CAS_19_23( {OUT_19_22[0], OUT_18_22[1], M[23], Q[13]}, OUT_19_23);
	wire [3:0] OUT_19_24;
	CAS CAS_19_24( {OUT_19_23[0], OUT_18_23[1], M[24], Q[13]}, OUT_19_24);
	wire [3:0] OUT_19_25;
	CAS CAS_19_25( {OUT_19_24[0], OUT_18_24[1], M[25], Q[13]}, OUT_19_25);
	wire [3:0] OUT_19_26;
	CAS CAS_19_26( {OUT_19_25[0], OUT_18_25[1], M[26], Q[13]}, OUT_19_26);
	wire [3:0] OUT_19_27;
	CAS CAS_19_27( {OUT_19_26[0], OUT_18_26[1], M[27], Q[13]}, OUT_19_27);
	wire [3:0] OUT_19_28;
	CAS CAS_19_28( {OUT_19_27[0], OUT_18_27[1], M[28], Q[13]}, OUT_19_28);
	wire [3:0] OUT_19_29;
	CAS CAS_19_29( {OUT_19_28[0], OUT_18_28[1], M[29], Q[13]}, OUT_19_29);
	wire [3:0] OUT_19_30;
	CAS CAS_19_30( {OUT_19_29[0], OUT_18_29[1], M[30], Q[13]}, OUT_19_30);
	wire [3:0] OUT_19_31;
	CAS CAS_19_31( {OUT_19_30[0], OUT_18_30[1], M[31], Q[13]}, OUT_19_31);
	assign Q[12] = OUT_19_31[0];

// Level - 21
	wire [3:0] OUT_20_0;
	CAS CAS_20_0( {Q[12], D[11], M[0], Q[12]}, OUT_20_0);
	wire [3:0] OUT_20_1;
	CAS CAS_20_1( {OUT_20_0[0], OUT_19_0[1], M[1], Q[12]}, OUT_20_1);
	wire [3:0] OUT_20_2;
	CAS CAS_20_2( {OUT_20_1[0], OUT_19_1[1], M[2], Q[12]}, OUT_20_2);
	wire [3:0] OUT_20_3;
	CAS CAS_20_3( {OUT_20_2[0], OUT_19_2[1], M[3], Q[12]}, OUT_20_3);
	wire [3:0] OUT_20_4;
	CAS CAS_20_4( {OUT_20_3[0], OUT_19_3[1], M[4], Q[12]}, OUT_20_4);
	wire [3:0] OUT_20_5;
	CAS CAS_20_5( {OUT_20_4[0], OUT_19_4[1], M[5], Q[12]}, OUT_20_5);
	wire [3:0] OUT_20_6;
	CAS CAS_20_6( {OUT_20_5[0], OUT_19_5[1], M[6], Q[12]}, OUT_20_6);
	wire [3:0] OUT_20_7;
	CAS CAS_20_7( {OUT_20_6[0], OUT_19_6[1], M[7], Q[12]}, OUT_20_7);
	wire [3:0] OUT_20_8;
	CAS CAS_20_8( {OUT_20_7[0], OUT_19_7[1], M[8], Q[12]}, OUT_20_8);
	wire [3:0] OUT_20_9;
	CAS CAS_20_9( {OUT_20_8[0], OUT_19_8[1], M[9], Q[12]}, OUT_20_9);
	wire [3:0] OUT_20_10;
	CAS CAS_20_10( {OUT_20_9[0], OUT_19_9[1], M[10], Q[12]}, OUT_20_10);
	wire [3:0] OUT_20_11;
	CAS CAS_20_11( {OUT_20_10[0], OUT_19_10[1], M[11], Q[12]}, OUT_20_11);
	wire [3:0] OUT_20_12;
	CAS CAS_20_12( {OUT_20_11[0], OUT_19_11[1], M[12], Q[12]}, OUT_20_12);
	wire [3:0] OUT_20_13;
	CAS CAS_20_13( {OUT_20_12[0], OUT_19_12[1], M[13], Q[12]}, OUT_20_13);
	wire [3:0] OUT_20_14;
	CAS CAS_20_14( {OUT_20_13[0], OUT_19_13[1], M[14], Q[12]}, OUT_20_14);
	wire [3:0] OUT_20_15;
	CAS CAS_20_15( {OUT_20_14[0], OUT_19_14[1], M[15], Q[12]}, OUT_20_15);
	wire [3:0] OUT_20_16;
	CAS CAS_20_16( {OUT_20_15[0], OUT_19_15[1], M[16], Q[12]}, OUT_20_16);
	wire [3:0] OUT_20_17;
	CAS CAS_20_17( {OUT_20_16[0], OUT_19_16[1], M[17], Q[12]}, OUT_20_17);
	wire [3:0] OUT_20_18;
	CAS CAS_20_18( {OUT_20_17[0], OUT_19_17[1], M[18], Q[12]}, OUT_20_18);
	wire [3:0] OUT_20_19;
	CAS CAS_20_19( {OUT_20_18[0], OUT_19_18[1], M[19], Q[12]}, OUT_20_19);
	wire [3:0] OUT_20_20;
	CAS CAS_20_20( {OUT_20_19[0], OUT_19_19[1], M[20], Q[12]}, OUT_20_20);
	wire [3:0] OUT_20_21;
	CAS CAS_20_21( {OUT_20_20[0], OUT_19_20[1], M[21], Q[12]}, OUT_20_21);
	wire [3:0] OUT_20_22;
	CAS CAS_20_22( {OUT_20_21[0], OUT_19_21[1], M[22], Q[12]}, OUT_20_22);
	wire [3:0] OUT_20_23;
	CAS CAS_20_23( {OUT_20_22[0], OUT_19_22[1], M[23], Q[12]}, OUT_20_23);
	wire [3:0] OUT_20_24;
	CAS CAS_20_24( {OUT_20_23[0], OUT_19_23[1], M[24], Q[12]}, OUT_20_24);
	wire [3:0] OUT_20_25;
	CAS CAS_20_25( {OUT_20_24[0], OUT_19_24[1], M[25], Q[12]}, OUT_20_25);
	wire [3:0] OUT_20_26;
	CAS CAS_20_26( {OUT_20_25[0], OUT_19_25[1], M[26], Q[12]}, OUT_20_26);
	wire [3:0] OUT_20_27;
	CAS CAS_20_27( {OUT_20_26[0], OUT_19_26[1], M[27], Q[12]}, OUT_20_27);
	wire [3:0] OUT_20_28;
	CAS CAS_20_28( {OUT_20_27[0], OUT_19_27[1], M[28], Q[12]}, OUT_20_28);
	wire [3:0] OUT_20_29;
	CAS CAS_20_29( {OUT_20_28[0], OUT_19_28[1], M[29], Q[12]}, OUT_20_29);
	wire [3:0] OUT_20_30;
	CAS CAS_20_30( {OUT_20_29[0], OUT_19_29[1], M[30], Q[12]}, OUT_20_30);
	wire [3:0] OUT_20_31;
	CAS CAS_20_31( {OUT_20_30[0], OUT_19_30[1], M[31], Q[12]}, OUT_20_31);
	assign Q[11] = OUT_20_31[0];

// Level - 22
	wire [3:0] OUT_21_0;
	CAS CAS_21_0( {Q[11], D[10], M[0], Q[11]}, OUT_21_0);
	wire [3:0] OUT_21_1;
	CAS CAS_21_1( {OUT_21_0[0], OUT_20_0[1], M[1], Q[11]}, OUT_21_1);
	wire [3:0] OUT_21_2;
	CAS CAS_21_2( {OUT_21_1[0], OUT_20_1[1], M[2], Q[11]}, OUT_21_2);
	wire [3:0] OUT_21_3;
	CAS CAS_21_3( {OUT_21_2[0], OUT_20_2[1], M[3], Q[11]}, OUT_21_3);
	wire [3:0] OUT_21_4;
	CAS CAS_21_4( {OUT_21_3[0], OUT_20_3[1], M[4], Q[11]}, OUT_21_4);
	wire [3:0] OUT_21_5;
	CAS CAS_21_5( {OUT_21_4[0], OUT_20_4[1], M[5], Q[11]}, OUT_21_5);
	wire [3:0] OUT_21_6;
	CAS CAS_21_6( {OUT_21_5[0], OUT_20_5[1], M[6], Q[11]}, OUT_21_6);
	wire [3:0] OUT_21_7;
	CAS CAS_21_7( {OUT_21_6[0], OUT_20_6[1], M[7], Q[11]}, OUT_21_7);
	wire [3:0] OUT_21_8;
	CAS CAS_21_8( {OUT_21_7[0], OUT_20_7[1], M[8], Q[11]}, OUT_21_8);
	wire [3:0] OUT_21_9;
	CAS CAS_21_9( {OUT_21_8[0], OUT_20_8[1], M[9], Q[11]}, OUT_21_9);
	wire [3:0] OUT_21_10;
	CAS CAS_21_10( {OUT_21_9[0], OUT_20_9[1], M[10], Q[11]}, OUT_21_10);
	wire [3:0] OUT_21_11;
	CAS CAS_21_11( {OUT_21_10[0], OUT_20_10[1], M[11], Q[11]}, OUT_21_11);
	wire [3:0] OUT_21_12;
	CAS CAS_21_12( {OUT_21_11[0], OUT_20_11[1], M[12], Q[11]}, OUT_21_12);
	wire [3:0] OUT_21_13;
	CAS CAS_21_13( {OUT_21_12[0], OUT_20_12[1], M[13], Q[11]}, OUT_21_13);
	wire [3:0] OUT_21_14;
	CAS CAS_21_14( {OUT_21_13[0], OUT_20_13[1], M[14], Q[11]}, OUT_21_14);
	wire [3:0] OUT_21_15;
	CAS CAS_21_15( {OUT_21_14[0], OUT_20_14[1], M[15], Q[11]}, OUT_21_15);
	wire [3:0] OUT_21_16;
	CAS CAS_21_16( {OUT_21_15[0], OUT_20_15[1], M[16], Q[11]}, OUT_21_16);
	wire [3:0] OUT_21_17;
	CAS CAS_21_17( {OUT_21_16[0], OUT_20_16[1], M[17], Q[11]}, OUT_21_17);
	wire [3:0] OUT_21_18;
	CAS CAS_21_18( {OUT_21_17[0], OUT_20_17[1], M[18], Q[11]}, OUT_21_18);
	wire [3:0] OUT_21_19;
	CAS CAS_21_19( {OUT_21_18[0], OUT_20_18[1], M[19], Q[11]}, OUT_21_19);
	wire [3:0] OUT_21_20;
	CAS CAS_21_20( {OUT_21_19[0], OUT_20_19[1], M[20], Q[11]}, OUT_21_20);
	wire [3:0] OUT_21_21;
	CAS CAS_21_21( {OUT_21_20[0], OUT_20_20[1], M[21], Q[11]}, OUT_21_21);
	wire [3:0] OUT_21_22;
	CAS CAS_21_22( {OUT_21_21[0], OUT_20_21[1], M[22], Q[11]}, OUT_21_22);
	wire [3:0] OUT_21_23;
	CAS CAS_21_23( {OUT_21_22[0], OUT_20_22[1], M[23], Q[11]}, OUT_21_23);
	wire [3:0] OUT_21_24;
	CAS CAS_21_24( {OUT_21_23[0], OUT_20_23[1], M[24], Q[11]}, OUT_21_24);
	wire [3:0] OUT_21_25;
	CAS CAS_21_25( {OUT_21_24[0], OUT_20_24[1], M[25], Q[11]}, OUT_21_25);
	wire [3:0] OUT_21_26;
	CAS CAS_21_26( {OUT_21_25[0], OUT_20_25[1], M[26], Q[11]}, OUT_21_26);
	wire [3:0] OUT_21_27;
	CAS CAS_21_27( {OUT_21_26[0], OUT_20_26[1], M[27], Q[11]}, OUT_21_27);
	wire [3:0] OUT_21_28;
	CAS CAS_21_28( {OUT_21_27[0], OUT_20_27[1], M[28], Q[11]}, OUT_21_28);
	wire [3:0] OUT_21_29;
	CAS CAS_21_29( {OUT_21_28[0], OUT_20_28[1], M[29], Q[11]}, OUT_21_29);
	wire [3:0] OUT_21_30;
	CAS CAS_21_30( {OUT_21_29[0], OUT_20_29[1], M[30], Q[11]}, OUT_21_30);
	wire [3:0] OUT_21_31;
	CAS CAS_21_31( {OUT_21_30[0], OUT_20_30[1], M[31], Q[11]}, OUT_21_31);
	assign Q[10] = OUT_21_31[0];

// Level - 23
	wire [3:0] OUT_22_0;
	CAS CAS_22_0( {Q[10], D[9], M[0], Q[10]}, OUT_22_0);
	wire [3:0] OUT_22_1;
	CAS CAS_22_1( {OUT_22_0[0], OUT_21_0[1], M[1], Q[10]}, OUT_22_1);
	wire [3:0] OUT_22_2;
	CAS CAS_22_2( {OUT_22_1[0], OUT_21_1[1], M[2], Q[10]}, OUT_22_2);
	wire [3:0] OUT_22_3;
	CAS CAS_22_3( {OUT_22_2[0], OUT_21_2[1], M[3], Q[10]}, OUT_22_3);
	wire [3:0] OUT_22_4;
	CAS CAS_22_4( {OUT_22_3[0], OUT_21_3[1], M[4], Q[10]}, OUT_22_4);
	wire [3:0] OUT_22_5;
	CAS CAS_22_5( {OUT_22_4[0], OUT_21_4[1], M[5], Q[10]}, OUT_22_5);
	wire [3:0] OUT_22_6;
	CAS CAS_22_6( {OUT_22_5[0], OUT_21_5[1], M[6], Q[10]}, OUT_22_6);
	wire [3:0] OUT_22_7;
	CAS CAS_22_7( {OUT_22_6[0], OUT_21_6[1], M[7], Q[10]}, OUT_22_7);
	wire [3:0] OUT_22_8;
	CAS CAS_22_8( {OUT_22_7[0], OUT_21_7[1], M[8], Q[10]}, OUT_22_8);
	wire [3:0] OUT_22_9;
	CAS CAS_22_9( {OUT_22_8[0], OUT_21_8[1], M[9], Q[10]}, OUT_22_9);
	wire [3:0] OUT_22_10;
	CAS CAS_22_10( {OUT_22_9[0], OUT_21_9[1], M[10], Q[10]}, OUT_22_10);
	wire [3:0] OUT_22_11;
	CAS CAS_22_11( {OUT_22_10[0], OUT_21_10[1], M[11], Q[10]}, OUT_22_11);
	wire [3:0] OUT_22_12;
	CAS CAS_22_12( {OUT_22_11[0], OUT_21_11[1], M[12], Q[10]}, OUT_22_12);
	wire [3:0] OUT_22_13;
	CAS CAS_22_13( {OUT_22_12[0], OUT_21_12[1], M[13], Q[10]}, OUT_22_13);
	wire [3:0] OUT_22_14;
	CAS CAS_22_14( {OUT_22_13[0], OUT_21_13[1], M[14], Q[10]}, OUT_22_14);
	wire [3:0] OUT_22_15;
	CAS CAS_22_15( {OUT_22_14[0], OUT_21_14[1], M[15], Q[10]}, OUT_22_15);
	wire [3:0] OUT_22_16;
	CAS CAS_22_16( {OUT_22_15[0], OUT_21_15[1], M[16], Q[10]}, OUT_22_16);
	wire [3:0] OUT_22_17;
	CAS CAS_22_17( {OUT_22_16[0], OUT_21_16[1], M[17], Q[10]}, OUT_22_17);
	wire [3:0] OUT_22_18;
	CAS CAS_22_18( {OUT_22_17[0], OUT_21_17[1], M[18], Q[10]}, OUT_22_18);
	wire [3:0] OUT_22_19;
	CAS CAS_22_19( {OUT_22_18[0], OUT_21_18[1], M[19], Q[10]}, OUT_22_19);
	wire [3:0] OUT_22_20;
	CAS CAS_22_20( {OUT_22_19[0], OUT_21_19[1], M[20], Q[10]}, OUT_22_20);
	wire [3:0] OUT_22_21;
	CAS CAS_22_21( {OUT_22_20[0], OUT_21_20[1], M[21], Q[10]}, OUT_22_21);
	wire [3:0] OUT_22_22;
	CAS CAS_22_22( {OUT_22_21[0], OUT_21_21[1], M[22], Q[10]}, OUT_22_22);
	wire [3:0] OUT_22_23;
	CAS CAS_22_23( {OUT_22_22[0], OUT_21_22[1], M[23], Q[10]}, OUT_22_23);
	wire [3:0] OUT_22_24;
	CAS CAS_22_24( {OUT_22_23[0], OUT_21_23[1], M[24], Q[10]}, OUT_22_24);
	wire [3:0] OUT_22_25;
	CAS CAS_22_25( {OUT_22_24[0], OUT_21_24[1], M[25], Q[10]}, OUT_22_25);
	wire [3:0] OUT_22_26;
	CAS CAS_22_26( {OUT_22_25[0], OUT_21_25[1], M[26], Q[10]}, OUT_22_26);
	wire [3:0] OUT_22_27;
	CAS CAS_22_27( {OUT_22_26[0], OUT_21_26[1], M[27], Q[10]}, OUT_22_27);
	wire [3:0] OUT_22_28;
	CAS CAS_22_28( {OUT_22_27[0], OUT_21_27[1], M[28], Q[10]}, OUT_22_28);
	wire [3:0] OUT_22_29;
	CAS CAS_22_29( {OUT_22_28[0], OUT_21_28[1], M[29], Q[10]}, OUT_22_29);
	wire [3:0] OUT_22_30;
	CAS CAS_22_30( {OUT_22_29[0], OUT_21_29[1], M[30], Q[10]}, OUT_22_30);
	wire [3:0] OUT_22_31;
	CAS CAS_22_31( {OUT_22_30[0], OUT_21_30[1], M[31], Q[10]}, OUT_22_31);
	assign Q[9] = OUT_22_31[0];

// Level - 24
	wire [3:0] OUT_23_0;
	CAS CAS_23_0( {Q[9], D[8], M[0], Q[9]}, OUT_23_0);
	wire [3:0] OUT_23_1;
	CAS CAS_23_1( {OUT_23_0[0], OUT_22_0[1], M[1], Q[9]}, OUT_23_1);
	wire [3:0] OUT_23_2;
	CAS CAS_23_2( {OUT_23_1[0], OUT_22_1[1], M[2], Q[9]}, OUT_23_2);
	wire [3:0] OUT_23_3;
	CAS CAS_23_3( {OUT_23_2[0], OUT_22_2[1], M[3], Q[9]}, OUT_23_3);
	wire [3:0] OUT_23_4;
	CAS CAS_23_4( {OUT_23_3[0], OUT_22_3[1], M[4], Q[9]}, OUT_23_4);
	wire [3:0] OUT_23_5;
	CAS CAS_23_5( {OUT_23_4[0], OUT_22_4[1], M[5], Q[9]}, OUT_23_5);
	wire [3:0] OUT_23_6;
	CAS CAS_23_6( {OUT_23_5[0], OUT_22_5[1], M[6], Q[9]}, OUT_23_6);
	wire [3:0] OUT_23_7;
	CAS CAS_23_7( {OUT_23_6[0], OUT_22_6[1], M[7], Q[9]}, OUT_23_7);
	wire [3:0] OUT_23_8;
	CAS CAS_23_8( {OUT_23_7[0], OUT_22_7[1], M[8], Q[9]}, OUT_23_8);
	wire [3:0] OUT_23_9;
	CAS CAS_23_9( {OUT_23_8[0], OUT_22_8[1], M[9], Q[9]}, OUT_23_9);
	wire [3:0] OUT_23_10;
	CAS CAS_23_10( {OUT_23_9[0], OUT_22_9[1], M[10], Q[9]}, OUT_23_10);
	wire [3:0] OUT_23_11;
	CAS CAS_23_11( {OUT_23_10[0], OUT_22_10[1], M[11], Q[9]}, OUT_23_11);
	wire [3:0] OUT_23_12;
	CAS CAS_23_12( {OUT_23_11[0], OUT_22_11[1], M[12], Q[9]}, OUT_23_12);
	wire [3:0] OUT_23_13;
	CAS CAS_23_13( {OUT_23_12[0], OUT_22_12[1], M[13], Q[9]}, OUT_23_13);
	wire [3:0] OUT_23_14;
	CAS CAS_23_14( {OUT_23_13[0], OUT_22_13[1], M[14], Q[9]}, OUT_23_14);
	wire [3:0] OUT_23_15;
	CAS CAS_23_15( {OUT_23_14[0], OUT_22_14[1], M[15], Q[9]}, OUT_23_15);
	wire [3:0] OUT_23_16;
	CAS CAS_23_16( {OUT_23_15[0], OUT_22_15[1], M[16], Q[9]}, OUT_23_16);
	wire [3:0] OUT_23_17;
	CAS CAS_23_17( {OUT_23_16[0], OUT_22_16[1], M[17], Q[9]}, OUT_23_17);
	wire [3:0] OUT_23_18;
	CAS CAS_23_18( {OUT_23_17[0], OUT_22_17[1], M[18], Q[9]}, OUT_23_18);
	wire [3:0] OUT_23_19;
	CAS CAS_23_19( {OUT_23_18[0], OUT_22_18[1], M[19], Q[9]}, OUT_23_19);
	wire [3:0] OUT_23_20;
	CAS CAS_23_20( {OUT_23_19[0], OUT_22_19[1], M[20], Q[9]}, OUT_23_20);
	wire [3:0] OUT_23_21;
	CAS CAS_23_21( {OUT_23_20[0], OUT_22_20[1], M[21], Q[9]}, OUT_23_21);
	wire [3:0] OUT_23_22;
	CAS CAS_23_22( {OUT_23_21[0], OUT_22_21[1], M[22], Q[9]}, OUT_23_22);
	wire [3:0] OUT_23_23;
	CAS CAS_23_23( {OUT_23_22[0], OUT_22_22[1], M[23], Q[9]}, OUT_23_23);
	wire [3:0] OUT_23_24;
	CAS CAS_23_24( {OUT_23_23[0], OUT_22_23[1], M[24], Q[9]}, OUT_23_24);
	wire [3:0] OUT_23_25;
	CAS CAS_23_25( {OUT_23_24[0], OUT_22_24[1], M[25], Q[9]}, OUT_23_25);
	wire [3:0] OUT_23_26;
	CAS CAS_23_26( {OUT_23_25[0], OUT_22_25[1], M[26], Q[9]}, OUT_23_26);
	wire [3:0] OUT_23_27;
	CAS CAS_23_27( {OUT_23_26[0], OUT_22_26[1], M[27], Q[9]}, OUT_23_27);
	wire [3:0] OUT_23_28;
	CAS CAS_23_28( {OUT_23_27[0], OUT_22_27[1], M[28], Q[9]}, OUT_23_28);
	wire [3:0] OUT_23_29;
	CAS CAS_23_29( {OUT_23_28[0], OUT_22_28[1], M[29], Q[9]}, OUT_23_29);
	wire [3:0] OUT_23_30;
	CAS CAS_23_30( {OUT_23_29[0], OUT_22_29[1], M[30], Q[9]}, OUT_23_30);
	wire [3:0] OUT_23_31;
	CAS CAS_23_31( {OUT_23_30[0], OUT_22_30[1], M[31], Q[9]}, OUT_23_31);
	assign Q[8] = OUT_23_31[0];

// Level - 25
	wire [3:0] OUT_24_0;
	CAS CAS_24_0( {Q[8], D[7], M[0], Q[8]}, OUT_24_0);
	wire [3:0] OUT_24_1;
	CAS CAS_24_1( {OUT_24_0[0], OUT_23_0[1], M[1], Q[8]}, OUT_24_1);
	wire [3:0] OUT_24_2;
	CAS CAS_24_2( {OUT_24_1[0], OUT_23_1[1], M[2], Q[8]}, OUT_24_2);
	wire [3:0] OUT_24_3;
	CAS CAS_24_3( {OUT_24_2[0], OUT_23_2[1], M[3], Q[8]}, OUT_24_3);
	wire [3:0] OUT_24_4;
	CAS CAS_24_4( {OUT_24_3[0], OUT_23_3[1], M[4], Q[8]}, OUT_24_4);
	wire [3:0] OUT_24_5;
	CAS CAS_24_5( {OUT_24_4[0], OUT_23_4[1], M[5], Q[8]}, OUT_24_5);
	wire [3:0] OUT_24_6;
	CAS CAS_24_6( {OUT_24_5[0], OUT_23_5[1], M[6], Q[8]}, OUT_24_6);
	wire [3:0] OUT_24_7;
	CAS CAS_24_7( {OUT_24_6[0], OUT_23_6[1], M[7], Q[8]}, OUT_24_7);
	wire [3:0] OUT_24_8;
	CAS CAS_24_8( {OUT_24_7[0], OUT_23_7[1], M[8], Q[8]}, OUT_24_8);
	wire [3:0] OUT_24_9;
	CAS CAS_24_9( {OUT_24_8[0], OUT_23_8[1], M[9], Q[8]}, OUT_24_9);
	wire [3:0] OUT_24_10;
	CAS CAS_24_10( {OUT_24_9[0], OUT_23_9[1], M[10], Q[8]}, OUT_24_10);
	wire [3:0] OUT_24_11;
	CAS CAS_24_11( {OUT_24_10[0], OUT_23_10[1], M[11], Q[8]}, OUT_24_11);
	wire [3:0] OUT_24_12;
	CAS CAS_24_12( {OUT_24_11[0], OUT_23_11[1], M[12], Q[8]}, OUT_24_12);
	wire [3:0] OUT_24_13;
	CAS CAS_24_13( {OUT_24_12[0], OUT_23_12[1], M[13], Q[8]}, OUT_24_13);
	wire [3:0] OUT_24_14;
	CAS CAS_24_14( {OUT_24_13[0], OUT_23_13[1], M[14], Q[8]}, OUT_24_14);
	wire [3:0] OUT_24_15;
	CAS CAS_24_15( {OUT_24_14[0], OUT_23_14[1], M[15], Q[8]}, OUT_24_15);
	wire [3:0] OUT_24_16;
	CAS CAS_24_16( {OUT_24_15[0], OUT_23_15[1], M[16], Q[8]}, OUT_24_16);
	wire [3:0] OUT_24_17;
	CAS CAS_24_17( {OUT_24_16[0], OUT_23_16[1], M[17], Q[8]}, OUT_24_17);
	wire [3:0] OUT_24_18;
	CAS CAS_24_18( {OUT_24_17[0], OUT_23_17[1], M[18], Q[8]}, OUT_24_18);
	wire [3:0] OUT_24_19;
	CAS CAS_24_19( {OUT_24_18[0], OUT_23_18[1], M[19], Q[8]}, OUT_24_19);
	wire [3:0] OUT_24_20;
	CAS CAS_24_20( {OUT_24_19[0], OUT_23_19[1], M[20], Q[8]}, OUT_24_20);
	wire [3:0] OUT_24_21;
	CAS CAS_24_21( {OUT_24_20[0], OUT_23_20[1], M[21], Q[8]}, OUT_24_21);
	wire [3:0] OUT_24_22;
	CAS CAS_24_22( {OUT_24_21[0], OUT_23_21[1], M[22], Q[8]}, OUT_24_22);
	wire [3:0] OUT_24_23;
	CAS CAS_24_23( {OUT_24_22[0], OUT_23_22[1], M[23], Q[8]}, OUT_24_23);
	wire [3:0] OUT_24_24;
	CAS CAS_24_24( {OUT_24_23[0], OUT_23_23[1], M[24], Q[8]}, OUT_24_24);
	wire [3:0] OUT_24_25;
	CAS CAS_24_25( {OUT_24_24[0], OUT_23_24[1], M[25], Q[8]}, OUT_24_25);
	wire [3:0] OUT_24_26;
	CAS CAS_24_26( {OUT_24_25[0], OUT_23_25[1], M[26], Q[8]}, OUT_24_26);
	wire [3:0] OUT_24_27;
	CAS CAS_24_27( {OUT_24_26[0], OUT_23_26[1], M[27], Q[8]}, OUT_24_27);
	wire [3:0] OUT_24_28;
	CAS CAS_24_28( {OUT_24_27[0], OUT_23_27[1], M[28], Q[8]}, OUT_24_28);
	wire [3:0] OUT_24_29;
	CAS CAS_24_29( {OUT_24_28[0], OUT_23_28[1], M[29], Q[8]}, OUT_24_29);
	wire [3:0] OUT_24_30;
	CAS CAS_24_30( {OUT_24_29[0], OUT_23_29[1], M[30], Q[8]}, OUT_24_30);
	wire [3:0] OUT_24_31;
	CAS CAS_24_31( {OUT_24_30[0], OUT_23_30[1], M[31], Q[8]}, OUT_24_31);
	assign Q[7] = OUT_24_31[0];

// Level - 26
	wire [3:0] OUT_25_0;
	CAS CAS_25_0( {Q[7], D[6], M[0], Q[7]}, OUT_25_0);
	wire [3:0] OUT_25_1;
	CAS CAS_25_1( {OUT_25_0[0], OUT_24_0[1], M[1], Q[7]}, OUT_25_1);
	wire [3:0] OUT_25_2;
	CAS CAS_25_2( {OUT_25_1[0], OUT_24_1[1], M[2], Q[7]}, OUT_25_2);
	wire [3:0] OUT_25_3;
	CAS CAS_25_3( {OUT_25_2[0], OUT_24_2[1], M[3], Q[7]}, OUT_25_3);
	wire [3:0] OUT_25_4;
	CAS CAS_25_4( {OUT_25_3[0], OUT_24_3[1], M[4], Q[7]}, OUT_25_4);
	wire [3:0] OUT_25_5;
	CAS CAS_25_5( {OUT_25_4[0], OUT_24_4[1], M[5], Q[7]}, OUT_25_5);
	wire [3:0] OUT_25_6;
	CAS CAS_25_6( {OUT_25_5[0], OUT_24_5[1], M[6], Q[7]}, OUT_25_6);
	wire [3:0] OUT_25_7;
	CAS CAS_25_7( {OUT_25_6[0], OUT_24_6[1], M[7], Q[7]}, OUT_25_7);
	wire [3:0] OUT_25_8;
	CAS CAS_25_8( {OUT_25_7[0], OUT_24_7[1], M[8], Q[7]}, OUT_25_8);
	wire [3:0] OUT_25_9;
	CAS CAS_25_9( {OUT_25_8[0], OUT_24_8[1], M[9], Q[7]}, OUT_25_9);
	wire [3:0] OUT_25_10;
	CAS CAS_25_10( {OUT_25_9[0], OUT_24_9[1], M[10], Q[7]}, OUT_25_10);
	wire [3:0] OUT_25_11;
	CAS CAS_25_11( {OUT_25_10[0], OUT_24_10[1], M[11], Q[7]}, OUT_25_11);
	wire [3:0] OUT_25_12;
	CAS CAS_25_12( {OUT_25_11[0], OUT_24_11[1], M[12], Q[7]}, OUT_25_12);
	wire [3:0] OUT_25_13;
	CAS CAS_25_13( {OUT_25_12[0], OUT_24_12[1], M[13], Q[7]}, OUT_25_13);
	wire [3:0] OUT_25_14;
	CAS CAS_25_14( {OUT_25_13[0], OUT_24_13[1], M[14], Q[7]}, OUT_25_14);
	wire [3:0] OUT_25_15;
	CAS CAS_25_15( {OUT_25_14[0], OUT_24_14[1], M[15], Q[7]}, OUT_25_15);
	wire [3:0] OUT_25_16;
	CAS CAS_25_16( {OUT_25_15[0], OUT_24_15[1], M[16], Q[7]}, OUT_25_16);
	wire [3:0] OUT_25_17;
	CAS CAS_25_17( {OUT_25_16[0], OUT_24_16[1], M[17], Q[7]}, OUT_25_17);
	wire [3:0] OUT_25_18;
	CAS CAS_25_18( {OUT_25_17[0], OUT_24_17[1], M[18], Q[7]}, OUT_25_18);
	wire [3:0] OUT_25_19;
	CAS CAS_25_19( {OUT_25_18[0], OUT_24_18[1], M[19], Q[7]}, OUT_25_19);
	wire [3:0] OUT_25_20;
	CAS CAS_25_20( {OUT_25_19[0], OUT_24_19[1], M[20], Q[7]}, OUT_25_20);
	wire [3:0] OUT_25_21;
	CAS CAS_25_21( {OUT_25_20[0], OUT_24_20[1], M[21], Q[7]}, OUT_25_21);
	wire [3:0] OUT_25_22;
	CAS CAS_25_22( {OUT_25_21[0], OUT_24_21[1], M[22], Q[7]}, OUT_25_22);
	wire [3:0] OUT_25_23;
	CAS CAS_25_23( {OUT_25_22[0], OUT_24_22[1], M[23], Q[7]}, OUT_25_23);
	wire [3:0] OUT_25_24;
	CAS CAS_25_24( {OUT_25_23[0], OUT_24_23[1], M[24], Q[7]}, OUT_25_24);
	wire [3:0] OUT_25_25;
	CAS CAS_25_25( {OUT_25_24[0], OUT_24_24[1], M[25], Q[7]}, OUT_25_25);
	wire [3:0] OUT_25_26;
	CAS CAS_25_26( {OUT_25_25[0], OUT_24_25[1], M[26], Q[7]}, OUT_25_26);
	wire [3:0] OUT_25_27;
	CAS CAS_25_27( {OUT_25_26[0], OUT_24_26[1], M[27], Q[7]}, OUT_25_27);
	wire [3:0] OUT_25_28;
	CAS CAS_25_28( {OUT_25_27[0], OUT_24_27[1], M[28], Q[7]}, OUT_25_28);
	wire [3:0] OUT_25_29;
	CAS CAS_25_29( {OUT_25_28[0], OUT_24_28[1], M[29], Q[7]}, OUT_25_29);
	wire [3:0] OUT_25_30;
	CAS CAS_25_30( {OUT_25_29[0], OUT_24_29[1], M[30], Q[7]}, OUT_25_30);
	wire [3:0] OUT_25_31;
	CAS CAS_25_31( {OUT_25_30[0], OUT_24_30[1], M[31], Q[7]}, OUT_25_31);
	assign Q[6] = OUT_25_31[0];

// Level - 27
	wire [3:0] OUT_26_0;
	CAS CAS_26_0( {Q[6], D[5], M[0], Q[6]}, OUT_26_0);
	wire [3:0] OUT_26_1;
	CAS CAS_26_1( {OUT_26_0[0], OUT_25_0[1], M[1], Q[6]}, OUT_26_1);
	wire [3:0] OUT_26_2;
	CAS CAS_26_2( {OUT_26_1[0], OUT_25_1[1], M[2], Q[6]}, OUT_26_2);
	wire [3:0] OUT_26_3;
	CAS CAS_26_3( {OUT_26_2[0], OUT_25_2[1], M[3], Q[6]}, OUT_26_3);
	wire [3:0] OUT_26_4;
	CAS CAS_26_4( {OUT_26_3[0], OUT_25_3[1], M[4], Q[6]}, OUT_26_4);
	wire [3:0] OUT_26_5;
	CAS CAS_26_5( {OUT_26_4[0], OUT_25_4[1], M[5], Q[6]}, OUT_26_5);
	wire [3:0] OUT_26_6;
	CAS CAS_26_6( {OUT_26_5[0], OUT_25_5[1], M[6], Q[6]}, OUT_26_6);
	wire [3:0] OUT_26_7;
	CAS CAS_26_7( {OUT_26_6[0], OUT_25_6[1], M[7], Q[6]}, OUT_26_7);
	wire [3:0] OUT_26_8;
	CAS CAS_26_8( {OUT_26_7[0], OUT_25_7[1], M[8], Q[6]}, OUT_26_8);
	wire [3:0] OUT_26_9;
	CAS CAS_26_9( {OUT_26_8[0], OUT_25_8[1], M[9], Q[6]}, OUT_26_9);
	wire [3:0] OUT_26_10;
	CAS CAS_26_10( {OUT_26_9[0], OUT_25_9[1], M[10], Q[6]}, OUT_26_10);
	wire [3:0] OUT_26_11;
	CAS CAS_26_11( {OUT_26_10[0], OUT_25_10[1], M[11], Q[6]}, OUT_26_11);
	wire [3:0] OUT_26_12;
	CAS CAS_26_12( {OUT_26_11[0], OUT_25_11[1], M[12], Q[6]}, OUT_26_12);
	wire [3:0] OUT_26_13;
	CAS CAS_26_13( {OUT_26_12[0], OUT_25_12[1], M[13], Q[6]}, OUT_26_13);
	wire [3:0] OUT_26_14;
	CAS CAS_26_14( {OUT_26_13[0], OUT_25_13[1], M[14], Q[6]}, OUT_26_14);
	wire [3:0] OUT_26_15;
	CAS CAS_26_15( {OUT_26_14[0], OUT_25_14[1], M[15], Q[6]}, OUT_26_15);
	wire [3:0] OUT_26_16;
	CAS CAS_26_16( {OUT_26_15[0], OUT_25_15[1], M[16], Q[6]}, OUT_26_16);
	wire [3:0] OUT_26_17;
	CAS CAS_26_17( {OUT_26_16[0], OUT_25_16[1], M[17], Q[6]}, OUT_26_17);
	wire [3:0] OUT_26_18;
	CAS CAS_26_18( {OUT_26_17[0], OUT_25_17[1], M[18], Q[6]}, OUT_26_18);
	wire [3:0] OUT_26_19;
	CAS CAS_26_19( {OUT_26_18[0], OUT_25_18[1], M[19], Q[6]}, OUT_26_19);
	wire [3:0] OUT_26_20;
	CAS CAS_26_20( {OUT_26_19[0], OUT_25_19[1], M[20], Q[6]}, OUT_26_20);
	wire [3:0] OUT_26_21;
	CAS CAS_26_21( {OUT_26_20[0], OUT_25_20[1], M[21], Q[6]}, OUT_26_21);
	wire [3:0] OUT_26_22;
	CAS CAS_26_22( {OUT_26_21[0], OUT_25_21[1], M[22], Q[6]}, OUT_26_22);
	wire [3:0] OUT_26_23;
	CAS CAS_26_23( {OUT_26_22[0], OUT_25_22[1], M[23], Q[6]}, OUT_26_23);
	wire [3:0] OUT_26_24;
	CAS CAS_26_24( {OUT_26_23[0], OUT_25_23[1], M[24], Q[6]}, OUT_26_24);
	wire [3:0] OUT_26_25;
	CAS CAS_26_25( {OUT_26_24[0], OUT_25_24[1], M[25], Q[6]}, OUT_26_25);
	wire [3:0] OUT_26_26;
	CAS CAS_26_26( {OUT_26_25[0], OUT_25_25[1], M[26], Q[6]}, OUT_26_26);
	wire [3:0] OUT_26_27;
	CAS CAS_26_27( {OUT_26_26[0], OUT_25_26[1], M[27], Q[6]}, OUT_26_27);
	wire [3:0] OUT_26_28;
	CAS CAS_26_28( {OUT_26_27[0], OUT_25_27[1], M[28], Q[6]}, OUT_26_28);
	wire [3:0] OUT_26_29;
	CAS CAS_26_29( {OUT_26_28[0], OUT_25_28[1], M[29], Q[6]}, OUT_26_29);
	wire [3:0] OUT_26_30;
	CAS CAS_26_30( {OUT_26_29[0], OUT_25_29[1], M[30], Q[6]}, OUT_26_30);
	wire [3:0] OUT_26_31;
	CAS CAS_26_31( {OUT_26_30[0], OUT_25_30[1], M[31], Q[6]}, OUT_26_31);
	assign Q[5] = OUT_26_31[0];

// Level - 28
	wire [3:0] OUT_27_0;
	CAS CAS_27_0( {Q[5], D[4], M[0], Q[5]}, OUT_27_0);
	wire [3:0] OUT_27_1;
	CAS CAS_27_1( {OUT_27_0[0], OUT_26_0[1], M[1], Q[5]}, OUT_27_1);
	wire [3:0] OUT_27_2;
	CAS CAS_27_2( {OUT_27_1[0], OUT_26_1[1], M[2], Q[5]}, OUT_27_2);
	wire [3:0] OUT_27_3;
	CAS CAS_27_3( {OUT_27_2[0], OUT_26_2[1], M[3], Q[5]}, OUT_27_3);
	wire [3:0] OUT_27_4;
	CAS CAS_27_4( {OUT_27_3[0], OUT_26_3[1], M[4], Q[5]}, OUT_27_4);
	wire [3:0] OUT_27_5;
	CAS CAS_27_5( {OUT_27_4[0], OUT_26_4[1], M[5], Q[5]}, OUT_27_5);
	wire [3:0] OUT_27_6;
	CAS CAS_27_6( {OUT_27_5[0], OUT_26_5[1], M[6], Q[5]}, OUT_27_6);
	wire [3:0] OUT_27_7;
	CAS CAS_27_7( {OUT_27_6[0], OUT_26_6[1], M[7], Q[5]}, OUT_27_7);
	wire [3:0] OUT_27_8;
	CAS CAS_27_8( {OUT_27_7[0], OUT_26_7[1], M[8], Q[5]}, OUT_27_8);
	wire [3:0] OUT_27_9;
	CAS CAS_27_9( {OUT_27_8[0], OUT_26_8[1], M[9], Q[5]}, OUT_27_9);
	wire [3:0] OUT_27_10;
	CAS CAS_27_10( {OUT_27_9[0], OUT_26_9[1], M[10], Q[5]}, OUT_27_10);
	wire [3:0] OUT_27_11;
	CAS CAS_27_11( {OUT_27_10[0], OUT_26_10[1], M[11], Q[5]}, OUT_27_11);
	wire [3:0] OUT_27_12;
	CAS CAS_27_12( {OUT_27_11[0], OUT_26_11[1], M[12], Q[5]}, OUT_27_12);
	wire [3:0] OUT_27_13;
	CAS CAS_27_13( {OUT_27_12[0], OUT_26_12[1], M[13], Q[5]}, OUT_27_13);
	wire [3:0] OUT_27_14;
	CAS CAS_27_14( {OUT_27_13[0], OUT_26_13[1], M[14], Q[5]}, OUT_27_14);
	wire [3:0] OUT_27_15;
	CAS CAS_27_15( {OUT_27_14[0], OUT_26_14[1], M[15], Q[5]}, OUT_27_15);
	wire [3:0] OUT_27_16;
	CAS CAS_27_16( {OUT_27_15[0], OUT_26_15[1], M[16], Q[5]}, OUT_27_16);
	wire [3:0] OUT_27_17;
	CAS CAS_27_17( {OUT_27_16[0], OUT_26_16[1], M[17], Q[5]}, OUT_27_17);
	wire [3:0] OUT_27_18;
	CAS CAS_27_18( {OUT_27_17[0], OUT_26_17[1], M[18], Q[5]}, OUT_27_18);
	wire [3:0] OUT_27_19;
	CAS CAS_27_19( {OUT_27_18[0], OUT_26_18[1], M[19], Q[5]}, OUT_27_19);
	wire [3:0] OUT_27_20;
	CAS CAS_27_20( {OUT_27_19[0], OUT_26_19[1], M[20], Q[5]}, OUT_27_20);
	wire [3:0] OUT_27_21;
	CAS CAS_27_21( {OUT_27_20[0], OUT_26_20[1], M[21], Q[5]}, OUT_27_21);
	wire [3:0] OUT_27_22;
	CAS CAS_27_22( {OUT_27_21[0], OUT_26_21[1], M[22], Q[5]}, OUT_27_22);
	wire [3:0] OUT_27_23;
	CAS CAS_27_23( {OUT_27_22[0], OUT_26_22[1], M[23], Q[5]}, OUT_27_23);
	wire [3:0] OUT_27_24;
	CAS CAS_27_24( {OUT_27_23[0], OUT_26_23[1], M[24], Q[5]}, OUT_27_24);
	wire [3:0] OUT_27_25;
	CAS CAS_27_25( {OUT_27_24[0], OUT_26_24[1], M[25], Q[5]}, OUT_27_25);
	wire [3:0] OUT_27_26;
	CAS CAS_27_26( {OUT_27_25[0], OUT_26_25[1], M[26], Q[5]}, OUT_27_26);
	wire [3:0] OUT_27_27;
	CAS CAS_27_27( {OUT_27_26[0], OUT_26_26[1], M[27], Q[5]}, OUT_27_27);
	wire [3:0] OUT_27_28;
	CAS CAS_27_28( {OUT_27_27[0], OUT_26_27[1], M[28], Q[5]}, OUT_27_28);
	wire [3:0] OUT_27_29;
	CAS CAS_27_29( {OUT_27_28[0], OUT_26_28[1], M[29], Q[5]}, OUT_27_29);
	wire [3:0] OUT_27_30;
	CAS CAS_27_30( {OUT_27_29[0], OUT_26_29[1], M[30], Q[5]}, OUT_27_30);
	wire [3:0] OUT_27_31;
	CAS CAS_27_31( {OUT_27_30[0], OUT_26_30[1], M[31], Q[5]}, OUT_27_31);
	assign Q[4] = OUT_27_31[0];

// Level - 29
	wire [3:0] OUT_28_0;
	CAS CAS_28_0( {Q[4], D[3], M[0], Q[4]}, OUT_28_0);
	wire [3:0] OUT_28_1;
	CAS CAS_28_1( {OUT_28_0[0], OUT_27_0[1], M[1], Q[4]}, OUT_28_1);
	wire [3:0] OUT_28_2;
	CAS CAS_28_2( {OUT_28_1[0], OUT_27_1[1], M[2], Q[4]}, OUT_28_2);
	wire [3:0] OUT_28_3;
	CAS CAS_28_3( {OUT_28_2[0], OUT_27_2[1], M[3], Q[4]}, OUT_28_3);
	wire [3:0] OUT_28_4;
	CAS CAS_28_4( {OUT_28_3[0], OUT_27_3[1], M[4], Q[4]}, OUT_28_4);
	wire [3:0] OUT_28_5;
	CAS CAS_28_5( {OUT_28_4[0], OUT_27_4[1], M[5], Q[4]}, OUT_28_5);
	wire [3:0] OUT_28_6;
	CAS CAS_28_6( {OUT_28_5[0], OUT_27_5[1], M[6], Q[4]}, OUT_28_6);
	wire [3:0] OUT_28_7;
	CAS CAS_28_7( {OUT_28_6[0], OUT_27_6[1], M[7], Q[4]}, OUT_28_7);
	wire [3:0] OUT_28_8;
	CAS CAS_28_8( {OUT_28_7[0], OUT_27_7[1], M[8], Q[4]}, OUT_28_8);
	wire [3:0] OUT_28_9;
	CAS CAS_28_9( {OUT_28_8[0], OUT_27_8[1], M[9], Q[4]}, OUT_28_9);
	wire [3:0] OUT_28_10;
	CAS CAS_28_10( {OUT_28_9[0], OUT_27_9[1], M[10], Q[4]}, OUT_28_10);
	wire [3:0] OUT_28_11;
	CAS CAS_28_11( {OUT_28_10[0], OUT_27_10[1], M[11], Q[4]}, OUT_28_11);
	wire [3:0] OUT_28_12;
	CAS CAS_28_12( {OUT_28_11[0], OUT_27_11[1], M[12], Q[4]}, OUT_28_12);
	wire [3:0] OUT_28_13;
	CAS CAS_28_13( {OUT_28_12[0], OUT_27_12[1], M[13], Q[4]}, OUT_28_13);
	wire [3:0] OUT_28_14;
	CAS CAS_28_14( {OUT_28_13[0], OUT_27_13[1], M[14], Q[4]}, OUT_28_14);
	wire [3:0] OUT_28_15;
	CAS CAS_28_15( {OUT_28_14[0], OUT_27_14[1], M[15], Q[4]}, OUT_28_15);
	wire [3:0] OUT_28_16;
	CAS CAS_28_16( {OUT_28_15[0], OUT_27_15[1], M[16], Q[4]}, OUT_28_16);
	wire [3:0] OUT_28_17;
	CAS CAS_28_17( {OUT_28_16[0], OUT_27_16[1], M[17], Q[4]}, OUT_28_17);
	wire [3:0] OUT_28_18;
	CAS CAS_28_18( {OUT_28_17[0], OUT_27_17[1], M[18], Q[4]}, OUT_28_18);
	wire [3:0] OUT_28_19;
	CAS CAS_28_19( {OUT_28_18[0], OUT_27_18[1], M[19], Q[4]}, OUT_28_19);
	wire [3:0] OUT_28_20;
	CAS CAS_28_20( {OUT_28_19[0], OUT_27_19[1], M[20], Q[4]}, OUT_28_20);
	wire [3:0] OUT_28_21;
	CAS CAS_28_21( {OUT_28_20[0], OUT_27_20[1], M[21], Q[4]}, OUT_28_21);
	wire [3:0] OUT_28_22;
	CAS CAS_28_22( {OUT_28_21[0], OUT_27_21[1], M[22], Q[4]}, OUT_28_22);
	wire [3:0] OUT_28_23;
	CAS CAS_28_23( {OUT_28_22[0], OUT_27_22[1], M[23], Q[4]}, OUT_28_23);
	wire [3:0] OUT_28_24;
	CAS CAS_28_24( {OUT_28_23[0], OUT_27_23[1], M[24], Q[4]}, OUT_28_24);
	wire [3:0] OUT_28_25;
	CAS CAS_28_25( {OUT_28_24[0], OUT_27_24[1], M[25], Q[4]}, OUT_28_25);
	wire [3:0] OUT_28_26;
	CAS CAS_28_26( {OUT_28_25[0], OUT_27_25[1], M[26], Q[4]}, OUT_28_26);
	wire [3:0] OUT_28_27;
	CAS CAS_28_27( {OUT_28_26[0], OUT_27_26[1], M[27], Q[4]}, OUT_28_27);
	wire [3:0] OUT_28_28;
	CAS CAS_28_28( {OUT_28_27[0], OUT_27_27[1], M[28], Q[4]}, OUT_28_28);
	wire [3:0] OUT_28_29;
	CAS CAS_28_29( {OUT_28_28[0], OUT_27_28[1], M[29], Q[4]}, OUT_28_29);
	wire [3:0] OUT_28_30;
	CAS CAS_28_30( {OUT_28_29[0], OUT_27_29[1], M[30], Q[4]}, OUT_28_30);
	wire [3:0] OUT_28_31;
	CAS CAS_28_31( {OUT_28_30[0], OUT_27_30[1], M[31], Q[4]}, OUT_28_31);
	assign Q[3] = OUT_28_31[0];

// Level - 30
	wire [3:0] OUT_29_0;
	CAS CAS_29_0( {Q[3], D[2], M[0], Q[3]}, OUT_29_0);
	wire [3:0] OUT_29_1;
	CAS CAS_29_1( {OUT_29_0[0], OUT_28_0[1], M[1], Q[3]}, OUT_29_1);
	wire [3:0] OUT_29_2;
	CAS CAS_29_2( {OUT_29_1[0], OUT_28_1[1], M[2], Q[3]}, OUT_29_2);
	wire [3:0] OUT_29_3;
	CAS CAS_29_3( {OUT_29_2[0], OUT_28_2[1], M[3], Q[3]}, OUT_29_3);
	wire [3:0] OUT_29_4;
	CAS CAS_29_4( {OUT_29_3[0], OUT_28_3[1], M[4], Q[3]}, OUT_29_4);
	wire [3:0] OUT_29_5;
	CAS CAS_29_5( {OUT_29_4[0], OUT_28_4[1], M[5], Q[3]}, OUT_29_5);
	wire [3:0] OUT_29_6;
	CAS CAS_29_6( {OUT_29_5[0], OUT_28_5[1], M[6], Q[3]}, OUT_29_6);
	wire [3:0] OUT_29_7;
	CAS CAS_29_7( {OUT_29_6[0], OUT_28_6[1], M[7], Q[3]}, OUT_29_7);
	wire [3:0] OUT_29_8;
	CAS CAS_29_8( {OUT_29_7[0], OUT_28_7[1], M[8], Q[3]}, OUT_29_8);
	wire [3:0] OUT_29_9;
	CAS CAS_29_9( {OUT_29_8[0], OUT_28_8[1], M[9], Q[3]}, OUT_29_9);
	wire [3:0] OUT_29_10;
	CAS CAS_29_10( {OUT_29_9[0], OUT_28_9[1], M[10], Q[3]}, OUT_29_10);
	wire [3:0] OUT_29_11;
	CAS CAS_29_11( {OUT_29_10[0], OUT_28_10[1], M[11], Q[3]}, OUT_29_11);
	wire [3:0] OUT_29_12;
	CAS CAS_29_12( {OUT_29_11[0], OUT_28_11[1], M[12], Q[3]}, OUT_29_12);
	wire [3:0] OUT_29_13;
	CAS CAS_29_13( {OUT_29_12[0], OUT_28_12[1], M[13], Q[3]}, OUT_29_13);
	wire [3:0] OUT_29_14;
	CAS CAS_29_14( {OUT_29_13[0], OUT_28_13[1], M[14], Q[3]}, OUT_29_14);
	wire [3:0] OUT_29_15;
	CAS CAS_29_15( {OUT_29_14[0], OUT_28_14[1], M[15], Q[3]}, OUT_29_15);
	wire [3:0] OUT_29_16;
	CAS CAS_29_16( {OUT_29_15[0], OUT_28_15[1], M[16], Q[3]}, OUT_29_16);
	wire [3:0] OUT_29_17;
	CAS CAS_29_17( {OUT_29_16[0], OUT_28_16[1], M[17], Q[3]}, OUT_29_17);
	wire [3:0] OUT_29_18;
	CAS CAS_29_18( {OUT_29_17[0], OUT_28_17[1], M[18], Q[3]}, OUT_29_18);
	wire [3:0] OUT_29_19;
	CAS CAS_29_19( {OUT_29_18[0], OUT_28_18[1], M[19], Q[3]}, OUT_29_19);
	wire [3:0] OUT_29_20;
	CAS CAS_29_20( {OUT_29_19[0], OUT_28_19[1], M[20], Q[3]}, OUT_29_20);
	wire [3:0] OUT_29_21;
	CAS CAS_29_21( {OUT_29_20[0], OUT_28_20[1], M[21], Q[3]}, OUT_29_21);
	wire [3:0] OUT_29_22;
	CAS CAS_29_22( {OUT_29_21[0], OUT_28_21[1], M[22], Q[3]}, OUT_29_22);
	wire [3:0] OUT_29_23;
	CAS CAS_29_23( {OUT_29_22[0], OUT_28_22[1], M[23], Q[3]}, OUT_29_23);
	wire [3:0] OUT_29_24;
	CAS CAS_29_24( {OUT_29_23[0], OUT_28_23[1], M[24], Q[3]}, OUT_29_24);
	wire [3:0] OUT_29_25;
	CAS CAS_29_25( {OUT_29_24[0], OUT_28_24[1], M[25], Q[3]}, OUT_29_25);
	wire [3:0] OUT_29_26;
	CAS CAS_29_26( {OUT_29_25[0], OUT_28_25[1], M[26], Q[3]}, OUT_29_26);
	wire [3:0] OUT_29_27;
	CAS CAS_29_27( {OUT_29_26[0], OUT_28_26[1], M[27], Q[3]}, OUT_29_27);
	wire [3:0] OUT_29_28;
	CAS CAS_29_28( {OUT_29_27[0], OUT_28_27[1], M[28], Q[3]}, OUT_29_28);
	wire [3:0] OUT_29_29;
	CAS CAS_29_29( {OUT_29_28[0], OUT_28_28[1], M[29], Q[3]}, OUT_29_29);
	wire [3:0] OUT_29_30;
	CAS CAS_29_30( {OUT_29_29[0], OUT_28_29[1], M[30], Q[3]}, OUT_29_30);
	wire [3:0] OUT_29_31;
	CAS CAS_29_31( {OUT_29_30[0], OUT_28_30[1], M[31], Q[3]}, OUT_29_31);
	assign Q[2] = OUT_29_31[0];

// Level - 31
	wire [3:0] OUT_30_0;
	CAS CAS_30_0( {Q[2], D[1], M[0], Q[2]}, OUT_30_0);
	wire [3:0] OUT_30_1;
	CAS CAS_30_1( {OUT_30_0[0], OUT_29_0[1], M[1], Q[2]}, OUT_30_1);
	wire [3:0] OUT_30_2;
	CAS CAS_30_2( {OUT_30_1[0], OUT_29_1[1], M[2], Q[2]}, OUT_30_2);
	wire [3:0] OUT_30_3;
	CAS CAS_30_3( {OUT_30_2[0], OUT_29_2[1], M[3], Q[2]}, OUT_30_3);
	wire [3:0] OUT_30_4;
	CAS CAS_30_4( {OUT_30_3[0], OUT_29_3[1], M[4], Q[2]}, OUT_30_4);
	wire [3:0] OUT_30_5;
	CAS CAS_30_5( {OUT_30_4[0], OUT_29_4[1], M[5], Q[2]}, OUT_30_5);
	wire [3:0] OUT_30_6;
	CAS CAS_30_6( {OUT_30_5[0], OUT_29_5[1], M[6], Q[2]}, OUT_30_6);
	wire [3:0] OUT_30_7;
	CAS CAS_30_7( {OUT_30_6[0], OUT_29_6[1], M[7], Q[2]}, OUT_30_7);
	wire [3:0] OUT_30_8;
	CAS CAS_30_8( {OUT_30_7[0], OUT_29_7[1], M[8], Q[2]}, OUT_30_8);
	wire [3:0] OUT_30_9;
	CAS CAS_30_9( {OUT_30_8[0], OUT_29_8[1], M[9], Q[2]}, OUT_30_9);
	wire [3:0] OUT_30_10;
	CAS CAS_30_10( {OUT_30_9[0], OUT_29_9[1], M[10], Q[2]}, OUT_30_10);
	wire [3:0] OUT_30_11;
	CAS CAS_30_11( {OUT_30_10[0], OUT_29_10[1], M[11], Q[2]}, OUT_30_11);
	wire [3:0] OUT_30_12;
	CAS CAS_30_12( {OUT_30_11[0], OUT_29_11[1], M[12], Q[2]}, OUT_30_12);
	wire [3:0] OUT_30_13;
	CAS CAS_30_13( {OUT_30_12[0], OUT_29_12[1], M[13], Q[2]}, OUT_30_13);
	wire [3:0] OUT_30_14;
	CAS CAS_30_14( {OUT_30_13[0], OUT_29_13[1], M[14], Q[2]}, OUT_30_14);
	wire [3:0] OUT_30_15;
	CAS CAS_30_15( {OUT_30_14[0], OUT_29_14[1], M[15], Q[2]}, OUT_30_15);
	wire [3:0] OUT_30_16;
	CAS CAS_30_16( {OUT_30_15[0], OUT_29_15[1], M[16], Q[2]}, OUT_30_16);
	wire [3:0] OUT_30_17;
	CAS CAS_30_17( {OUT_30_16[0], OUT_29_16[1], M[17], Q[2]}, OUT_30_17);
	wire [3:0] OUT_30_18;
	CAS CAS_30_18( {OUT_30_17[0], OUT_29_17[1], M[18], Q[2]}, OUT_30_18);
	wire [3:0] OUT_30_19;
	CAS CAS_30_19( {OUT_30_18[0], OUT_29_18[1], M[19], Q[2]}, OUT_30_19);
	wire [3:0] OUT_30_20;
	CAS CAS_30_20( {OUT_30_19[0], OUT_29_19[1], M[20], Q[2]}, OUT_30_20);
	wire [3:0] OUT_30_21;
	CAS CAS_30_21( {OUT_30_20[0], OUT_29_20[1], M[21], Q[2]}, OUT_30_21);
	wire [3:0] OUT_30_22;
	CAS CAS_30_22( {OUT_30_21[0], OUT_29_21[1], M[22], Q[2]}, OUT_30_22);
	wire [3:0] OUT_30_23;
	CAS CAS_30_23( {OUT_30_22[0], OUT_29_22[1], M[23], Q[2]}, OUT_30_23);
	wire [3:0] OUT_30_24;
	CAS CAS_30_24( {OUT_30_23[0], OUT_29_23[1], M[24], Q[2]}, OUT_30_24);
	wire [3:0] OUT_30_25;
	CAS CAS_30_25( {OUT_30_24[0], OUT_29_24[1], M[25], Q[2]}, OUT_30_25);
	wire [3:0] OUT_30_26;
	CAS CAS_30_26( {OUT_30_25[0], OUT_29_25[1], M[26], Q[2]}, OUT_30_26);
	wire [3:0] OUT_30_27;
	CAS CAS_30_27( {OUT_30_26[0], OUT_29_26[1], M[27], Q[2]}, OUT_30_27);
	wire [3:0] OUT_30_28;
	CAS CAS_30_28( {OUT_30_27[0], OUT_29_27[1], M[28], Q[2]}, OUT_30_28);
	wire [3:0] OUT_30_29;
	CAS CAS_30_29( {OUT_30_28[0], OUT_29_28[1], M[29], Q[2]}, OUT_30_29);
	wire [3:0] OUT_30_30;
	CAS CAS_30_30( {OUT_30_29[0], OUT_29_29[1], M[30], Q[2]}, OUT_30_30);
	wire [3:0] OUT_30_31;
	CAS CAS_30_31( {OUT_30_30[0], OUT_29_30[1], M[31], Q[2]}, OUT_30_31);
	assign Q[1] = OUT_30_31[0];

// Level - 32
	wire [3:0] OUT_31_0;
	CAS CAS_31_0( {Q[1], D[0], M[0], Q[1]}, OUT_31_0);
	wire [3:0] OUT_31_1;
	CAS CAS_31_1( {OUT_31_0[0], OUT_30_0[1], M[1], Q[1]}, OUT_31_1);
	wire [3:0] OUT_31_2;
	CAS CAS_31_2( {OUT_31_1[0], OUT_30_1[1], M[2], Q[1]}, OUT_31_2);
	wire [3:0] OUT_31_3;
	CAS CAS_31_3( {OUT_31_2[0], OUT_30_2[1], M[3], Q[1]}, OUT_31_3);
	wire [3:0] OUT_31_4;
	CAS CAS_31_4( {OUT_31_3[0], OUT_30_3[1], M[4], Q[1]}, OUT_31_4);
	wire [3:0] OUT_31_5;
	CAS CAS_31_5( {OUT_31_4[0], OUT_30_4[1], M[5], Q[1]}, OUT_31_5);
	wire [3:0] OUT_31_6;
	CAS CAS_31_6( {OUT_31_5[0], OUT_30_5[1], M[6], Q[1]}, OUT_31_6);
	wire [3:0] OUT_31_7;
	CAS CAS_31_7( {OUT_31_6[0], OUT_30_6[1], M[7], Q[1]}, OUT_31_7);
	wire [3:0] OUT_31_8;
	CAS CAS_31_8( {OUT_31_7[0], OUT_30_7[1], M[8], Q[1]}, OUT_31_8);
	wire [3:0] OUT_31_9;
	CAS CAS_31_9( {OUT_31_8[0], OUT_30_8[1], M[9], Q[1]}, OUT_31_9);
	wire [3:0] OUT_31_10;
	CAS CAS_31_10( {OUT_31_9[0], OUT_30_9[1], M[10], Q[1]}, OUT_31_10);
	wire [3:0] OUT_31_11;
	CAS CAS_31_11( {OUT_31_10[0], OUT_30_10[1], M[11], Q[1]}, OUT_31_11);
	wire [3:0] OUT_31_12;
	CAS CAS_31_12( {OUT_31_11[0], OUT_30_11[1], M[12], Q[1]}, OUT_31_12);
	wire [3:0] OUT_31_13;
	CAS CAS_31_13( {OUT_31_12[0], OUT_30_12[1], M[13], Q[1]}, OUT_31_13);
	wire [3:0] OUT_31_14;
	CAS CAS_31_14( {OUT_31_13[0], OUT_30_13[1], M[14], Q[1]}, OUT_31_14);
	wire [3:0] OUT_31_15;
	CAS CAS_31_15( {OUT_31_14[0], OUT_30_14[1], M[15], Q[1]}, OUT_31_15);
	wire [3:0] OUT_31_16;
	CAS CAS_31_16( {OUT_31_15[0], OUT_30_15[1], M[16], Q[1]}, OUT_31_16);
	wire [3:0] OUT_31_17;
	CAS CAS_31_17( {OUT_31_16[0], OUT_30_16[1], M[17], Q[1]}, OUT_31_17);
	wire [3:0] OUT_31_18;
	CAS CAS_31_18( {OUT_31_17[0], OUT_30_17[1], M[18], Q[1]}, OUT_31_18);
	wire [3:0] OUT_31_19;
	CAS CAS_31_19( {OUT_31_18[0], OUT_30_18[1], M[19], Q[1]}, OUT_31_19);
	wire [3:0] OUT_31_20;
	CAS CAS_31_20( {OUT_31_19[0], OUT_30_19[1], M[20], Q[1]}, OUT_31_20);
	wire [3:0] OUT_31_21;
	CAS CAS_31_21( {OUT_31_20[0], OUT_30_20[1], M[21], Q[1]}, OUT_31_21);
	wire [3:0] OUT_31_22;
	CAS CAS_31_22( {OUT_31_21[0], OUT_30_21[1], M[22], Q[1]}, OUT_31_22);
	wire [3:0] OUT_31_23;
	CAS CAS_31_23( {OUT_31_22[0], OUT_30_22[1], M[23], Q[1]}, OUT_31_23);
	wire [3:0] OUT_31_24;
	CAS CAS_31_24( {OUT_31_23[0], OUT_30_23[1], M[24], Q[1]}, OUT_31_24);
	wire [3:0] OUT_31_25;
	CAS CAS_31_25( {OUT_31_24[0], OUT_30_24[1], M[25], Q[1]}, OUT_31_25);
	wire [3:0] OUT_31_26;
	CAS CAS_31_26( {OUT_31_25[0], OUT_30_25[1], M[26], Q[1]}, OUT_31_26);
	wire [3:0] OUT_31_27;
	CAS CAS_31_27( {OUT_31_26[0], OUT_30_26[1], M[27], Q[1]}, OUT_31_27);
	wire [3:0] OUT_31_28;
	CAS CAS_31_28( {OUT_31_27[0], OUT_30_27[1], M[28], Q[1]}, OUT_31_28);
	wire [3:0] OUT_31_29;
	CAS CAS_31_29( {OUT_31_28[0], OUT_30_28[1], M[29], Q[1]}, OUT_31_29);
	wire [3:0] OUT_31_30;
	CAS CAS_31_30( {OUT_31_29[0], OUT_30_29[1], M[30], Q[1]}, OUT_31_30);
	wire [3:0] OUT_31_31;
	CAS CAS_31_31( {OUT_31_30[0], OUT_30_30[1], M[31], Q[1]}, OUT_31_31);
	assign Q[0] = OUT_31_31[0];

// Remainder Correction
	wire C_0 = 1'b0;
	assign R[0] = OUT_31_0[1] ^ ( M[0] & OUT_31_31[1]) ^ C_0;

	wire C_1 = (OUT_31_0[1] & ( M[0] & OUT_31_31[1])) | (C_0 & (OUT_31_0[1] ^( M[0] & OUT_31_31[1])));
        assign R[1] = OUT_31_1[1] ^ ( M[1] & OUT_31_31[1]) ^ C_1;

        wire C_2 = (OUT_31_1[1] & ( M[1] & OUT_31_31[1])) | (C_1 & (OUT_31_1[1] ^( M[1] & OUT_31_31[1])));
        assign R[2] = OUT_31_2[1] ^ ( M[2] & OUT_31_31[1]) ^ C_2;

wire C_3 = (OUT_31_2[1] & ( M[2] & OUT_31_31[1])) | (C_2 & (OUT_31_2[1] ^( M[2] & OUT_31_31[1])));
	assign R[3] = OUT_31_3[1] ^ ( M[3] & OUT_31_31[1]) ^ C_3;

	wire C_4 = (OUT_31_3[1] & ( M[3] & OUT_31_31[1])) | (C_3 & (OUT_31_3[1] ^( M[3] & OUT_31_31[1])));
	assign R[4] = OUT_31_4[1] ^ ( M[4] & OUT_31_31[1]) ^ C_4;

	wire C_5 = (OUT_31_4[1] & ( M[4] & OUT_31_31[1])) | (C_4 & (OUT_31_4[1] ^( M[4] & OUT_31_31[1])));
	assign R[5] = OUT_31_5[1] ^ ( M[5] & OUT_31_31[1]) ^ C_5;

	wire C_6 = (OUT_31_5[1] & ( M[5] & OUT_31_31[1])) | (C_5 & (OUT_31_5[1] ^( M[5] & OUT_31_31[1])));
	assign R[6] = OUT_31_6[1] ^ ( M[6] & OUT_31_31[1]) ^ C_6;

	wire C_7 = (OUT_31_6[1] & ( M[6] & OUT_31_31[1])) | (C_6 & (OUT_31_6[1] ^( M[6] & OUT_31_31[1])));
	assign R[7] = OUT_31_7[1] ^ ( M[7] & OUT_31_31[1]) ^ C_7;

	wire C_8 = (OUT_31_7[1] & ( M[7] & OUT_31_31[1])) | (C_7 & (OUT_31_7[1] ^( M[7] & OUT_31_31[1])));
	assign R[8] = OUT_31_8[1] ^ ( M[8] & OUT_31_31[1]) ^ C_8;

	wire C_9 = (OUT_31_8[1] & ( M[8] & OUT_31_31[1])) | (C_8 & (OUT_31_8[1] ^( M[8] & OUT_31_31[1])));
	assign R[9] = OUT_31_9[1] ^ ( M[9] & OUT_31_31[1]) ^ C_9;

	wire C_10 = (OUT_31_9[1] & ( M[9] & OUT_31_31[1])) | (C_9 & (OUT_31_9[1] ^( M[9] & OUT_31_31[1])));
	assign R[10] = OUT_31_10[1] ^ ( M[10] & OUT_31_31[1]) ^ C_10;

	wire C_11 = (OUT_31_10[1] & ( M[10] & OUT_31_31[1])) | (C_10 & (OUT_31_10[1] ^( M[10] & OUT_31_31[1])));
	assign R[11] = OUT_31_11[1] ^ ( M[11] & OUT_31_31[1]) ^ C_11;

	wire C_12 = (OUT_31_11[1] & ( M[11] & OUT_31_31[1])) | (C_11 & (OUT_31_11[1] ^( M[11] & OUT_31_31[1])));
	assign R[12] = OUT_31_12[1] ^ ( M[12] & OUT_31_31[1]) ^ C_12;

	wire C_13 = (OUT_31_12[1] & ( M[12] & OUT_31_31[1])) | (C_12 & (OUT_31_12[1] ^( M[12] & OUT_31_31[1])));
	assign R[13] = OUT_31_13[1] ^ ( M[13] & OUT_31_31[1]) ^ C_13;

	wire C_14 = (OUT_31_13[1] & ( M[13] & OUT_31_31[1])) | (C_13 & (OUT_31_13[1] ^( M[13] & OUT_31_31[1])));
	assign R[14] = OUT_31_14[1] ^ ( M[14] & OUT_31_31[1]) ^ C_14;

	wire C_15 = (OUT_31_14[1] & ( M[14] & OUT_31_31[1])) | (C_14 & (OUT_31_14[1] ^( M[14] & OUT_31_31[1])));
	assign R[15] = OUT_31_15[1] ^ ( M[15] & OUT_31_31[1]) ^ C_15;

	wire C_16 = (OUT_31_15[1] & ( M[15] & OUT_31_31[1])) | (C_15 & (OUT_31_15[1] ^( M[15] & OUT_31_31[1])));
	assign R[16] = OUT_31_16[1] ^ ( M[16] & OUT_31_31[1]) ^ C_16;

	wire C_17 = (OUT_31_16[1] & ( M[16] & OUT_31_31[1])) | (C_16 & (OUT_31_16[1] ^( M[16] & OUT_31_31[1])));
	assign R[17] = OUT_31_17[1] ^ ( M[17] & OUT_31_31[1]) ^ C_17;

	wire C_18 = (OUT_31_17[1] & ( M[17] & OUT_31_31[1])) | (C_17 & (OUT_31_17[1] ^( M[17] & OUT_31_31[1])));
	assign R[18] = OUT_31_18[1] ^ ( M[18] & OUT_31_31[1]) ^ C_18;

	wire C_19 = (OUT_31_18[1] & ( M[18] & OUT_31_31[1])) | (C_18 & (OUT_31_18[1] ^( M[18] & OUT_31_31[1])));
	assign R[19] = OUT_31_19[1] ^ ( M[19] & OUT_31_31[1]) ^ C_19;

	wire C_20 = (OUT_31_19[1] & ( M[19] & OUT_31_31[1])) | (C_19 & (OUT_31_19[1] ^( M[19] & OUT_31_31[1])));
	assign R[20] = OUT_31_20[1] ^ ( M[20] & OUT_31_31[1]) ^ C_20;

	wire C_21 = (OUT_31_20[1] & ( M[20] & OUT_31_31[1])) | (C_20 & (OUT_31_20[1] ^( M[20] & OUT_31_31[1])));
	assign R[21] = OUT_31_21[1] ^ ( M[21] & OUT_31_31[1]) ^ C_21;

	wire C_22 = (OUT_31_21[1] & ( M[21] & OUT_31_31[1])) | (C_21 & (OUT_31_21[1] ^( M[21] & OUT_31_31[1])));
	assign R[22] = OUT_31_22[1] ^ ( M[22] & OUT_31_31[1]) ^ C_22;

	wire C_23 = (OUT_31_22[1] & ( M[22] & OUT_31_31[1])) | (C_22 & (OUT_31_22[1] ^( M[22] & OUT_31_31[1])));
	assign R[23] = OUT_31_23[1] ^ ( M[23] & OUT_31_31[1]) ^ C_23;

	wire C_24 = (OUT_31_23[1] & ( M[23] & OUT_31_31[1])) | (C_23 & (OUT_31_23[1] ^( M[23] & OUT_31_31[1])));
	assign R[24] = OUT_31_24[1] ^ ( M[24] & OUT_31_31[1]) ^ C_24;

	wire C_25 = (OUT_31_24[1] & ( M[24] & OUT_31_31[1])) | (C_24 & (OUT_31_24[1] ^( M[24] & OUT_31_31[1])));
	assign R[25] = OUT_31_25[1] ^ ( M[25] & OUT_31_31[1]) ^ C_25;

	wire C_26 = (OUT_31_25[1] & ( M[25] & OUT_31_31[1])) | (C_25 & (OUT_31_25[1] ^( M[25] & OUT_31_31[1])));
	assign R[26] = OUT_31_26[1] ^ ( M[26] & OUT_31_31[1]) ^ C_26;

	wire C_27 = (OUT_31_26[1] & ( M[26] & OUT_31_31[1])) | (C_26 & (OUT_31_26[1] ^( M[26] & OUT_31_31[1])));
	assign R[27] = OUT_31_27[1] ^ ( M[27] & OUT_31_31[1]) ^ C_27;

	wire C_28 = (OUT_31_27[1] & ( M[27] & OUT_31_31[1])) | (C_27 & (OUT_31_27[1] ^( M[27] & OUT_31_31[1])));
	assign R[28] = OUT_31_28[1] ^ ( M[28] & OUT_31_31[1]) ^ C_28;

	wire C_29 = (OUT_31_28[1] & ( M[28] & OUT_31_31[1])) | (C_28 & (OUT_31_28[1] ^( M[28] & OUT_31_31[1])));
	assign R[29] = OUT_31_29[1] ^ ( M[29] & OUT_31_31[1]) ^ C_29;

	wire C_30 = (OUT_31_29[1] & ( M[29] & OUT_31_31[1])) | (C_29 & (OUT_31_29[1] ^( M[29] & OUT_31_31[1])));
	assign R[30] = OUT_31_30[1] ^ ( M[30] & OUT_31_31[1]) ^ C_30;

	wire C_31 = (OUT_31_30[1] & ( M[30] & OUT_31_31[1])) | (C_30 & (OUT_31_30[1] ^( M[30] & OUT_31_31[1])));
	assign R[31] = OUT_31_31[1] ^ ( M[31] & OUT_31_31[1]) ^ C_31;

endmodule

